* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 2
.param
+ sky130_fd_pr__special_nfet_01v8__toxe_mult = 1.0
+ sky130_fd_pr__special_nfet_01v8__rshn_mult = 1.0
+ sky130_fd_pr__special_nfet_01v8__overlap_mult = 0.9642
+ sky130_fd_pr__special_nfet_01v8__lint_diff = 0.0
+ sky130_fd_pr__special_nfet_01v8__wint_diff = 0.0
+ sky130_fd_pr__special_nfet_01v8__dlc_diff = -.61491e-9
+ sky130_fd_pr__special_nfet_01v8__dwc_diff = 0.0
*
* sky130_fd_pr__special_nfet_01v8, Bin 000, W = 0.36, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_01v8__ub_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vsat_diff_0 = 2522.7
+ sky130_fd_pr__special_nfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vth0_diff_0 = 0.042691
+ sky130_fd_pr__special_nfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__u0_diff_0 = 0.0031326
+ sky130_fd_pr__special_nfet_01v8__nfactor_diff_0 = 0.93967
+ sky130_fd_pr__special_nfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__k2_diff_0 = -0.011632
+ sky130_fd_pr__special_nfet_01v8__ua_diff_0 = 0.0
*
* sky130_fd_pr__special_nfet_01v8, Bin 001, W = 0.39, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_01v8__ua_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__ub_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vsat_diff_1 = 1928.2
+ sky130_fd_pr__special_nfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vth0_diff_1 = 0.032658
+ sky130_fd_pr__special_nfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b0_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__voff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__u0_diff_1 = 0.0029052
+ sky130_fd_pr__special_nfet_01v8__nfactor_diff_1 = 0.83163
+ sky130_fd_pr__special_nfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__ags_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__k2_diff_1 = -0.009063
*
.include "sky130_fd_pr__special_nfet_01v8.pm3.spice"
