* Copyright 2022 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SKY130 Device models.
*----------------------------------------------------------
* This file includes all legacy discrete models from the
* original skywater-pdk that are not included in the set
* of continuous models.
*
* This file is used for monte carlo process simulations.
* For corner and mismatch simulations, use "all.spice".
*----------------------------------------------------------
* The scale option forces all netlists to provide distance
* units in microns (e.g., 1 micron width is W=1, not W=1u).
* The first scale option is used by ngspice, the second by
* Xyce.  Each tool ignores the other's syntax.
*----------------------------------------------------------
.option scale=1.0u
.options parser scale=1.0u

.include "invariant.spice"

*----------------------------------------------------------
* Derivative Parameters:
*----------------------------------------------------------
.param
+ cnwvc2_cdepmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc2_cintmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc2_dlc = '-2.50000e-03*cnwvc'
+ cnwvc2_dld = '-1.50000e-04*cnwvc'
+ cnwvc2_dwc = '-5.00000e-03*cnwvc'
+ cnwvc2_tox = '1.32732e-02*cnwvc*cnwvc+5.84020e-01*cnwvc+4.24742e+01'
+ cnwvc2_vt1 = '1.85000e-02*cnwvc+2.00000e-01'
+ cnwvc2_vt2 = '1.85000e-02*cnwvc+3.30000e-01'
+ cnwvc2_vtr = '1.85000e-02*cnwvc+1.40000e-01'
+ cnwvc_cdepmult = '-2.50000e-02*cnwvc+1.00000e+00'
+ cnwvc_cintmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc_dlc = '-2.50000e-03*poly_cd'
+ cnwvc_dld = '-2.00000e-04*cnwvc'
+ cnwvc_dwc = '-5.00000e-03*cnwvc'
+ cnwvc_tox = '1.59937e-02*cnwvc*cnwvc+5.75774e-01*cnwvc+4.26499e+01'
+ cnwvc_vt1 = '2.80000e-02*lvp_threshold+3.33300e-01'
+ cnwvc_vt2 = '2.80000e-02*lvp_threshold+2.38095e-01'
+ cnwvc_vtr = '2.80000e-02*lvp_threshold+1.60000e-01'
+ c0m4m3_vpp = '9.09375e-03*ic_cap*ic_cap+8.53750e-02*ic_cap+1.00000e+00'
+ c0m5m3_vpp = '5.28125e-03*ic_cap*ic_cap+7.03750e-02*ic_cap+1.00000e+00'
+ c0m5m4_vpp = '9.09375e-03*ic_cap*ic_cap+8.53750e-02*ic_cap+1.00000e+00'
+ c0m5m4_vpp0p4shield = '5.14350e-02*ic_cap*ic_cap+3.04590e-01*ic_cap+1.00000e+00'
+ c1m4m3_vpp = '5.78125e-03*ic_cap*ic_cap+8.16250e-02*ic_cap+1.00000e+00'
+ c1m5m3_vpp = '8.43750e-03*ic_cap*ic_cap+9.02500e-02*ic_cap+1.00000e+00'
+ c1m5m4_vpp = '5.78125e-03*ic_cap*ic_cap+8.16250e-02*ic_cap+1.00000e+00'
+ c1m5m4_vpp0p4shield = '8.44188e-03*ic_cap*ic_cap+9.22675e-02*ic_cap+1.00000e+00'
+ cvpp2_nhvnative10x4_cor = '-6.25000e-05*ic_cap*ic_cap+-3.42500e-02*ic_cap+1.00000e+00'
+ cvpp2_nhvnative10x4_sub = '1.10250e-16*ic_cap*ic_cap+-1.42900e-15*ic_cap+4.82000e-15'
+ cvpp2_phv5x4_cor = '-6.25000e-05*ic_cap*ic_cap+-3.42500e-02*ic_cap+1.00000e+00'
+ cvpp2_phv5x4_sub = '1.10250e-16*ic_cap*ic_cap+-1.42900e-15*ic_cap+4.82000e-15'
+ cvpp3_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp4_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp5_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp_cor = '-6.25000e-05*ic_cap*ic_cap+3.42500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = '-2.50000e-06*hvp_diode*hvp_diode+1.81850e-02*hvp_diode+1.00500e+00'
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__nfet_05v0_nvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_20v0__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_20v0_nvt_iso__hvvsat_mult = '2.48544e-02*hvn_saturation*hvn_saturation+-5.96505e-02*hvn_saturation+1.00000e-18'
+ sky130_fd_pr__nfet_20v0_nvt_iso__rdrift_mult = '2.07703e-02*nfet_20v0_nvt_iso*nfet_20v0_nvt_iso+1.69501e-01*nfet_20v0_nvt_iso+8.20770e-01'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vth0_diff = '2.00325e-04*hvntvn_threshold*hvntvn_threshold+3.47038e-02*hvntvn_threshold+4.46980e-03'
+ sky130_fd_pr__special_nfet_pass_flash__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_pass_flash__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_flash__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1 = '-1.06270e-02*lvn_subvt*lvn_subvt+1.13538e-02*lvn_subvt+3.82270e-02'
+ sky130_fd_pr__special_nfet_pass_flash__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0 = '-7.91375e-03*lvn_subvt*lvn_subvt+3.16550e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1 = '1.41651e-02*lvn_subvt*lvn_subvt+8.47347e-02*lvn_subvt+1.41380e-01'
+ sky130_fd_pr__special_nfet_pass_flash__overlap_mult = '1.18750e-04*lvtox*lvtox+2.44075e-02*lvtox+8.98050e-01'
+ sky130_fd_pr__special_nfet_pass_flash__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_pass_flash__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_0 = '-1.24384e-05*lvn_mobility*lvn_mobility+8.14504e-04*lvn_mobility+2.75840e-03'
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_1 = '-1.68563e-04*lvn_mobility*lvn_mobility+1.84207e-03*lvn_mobility+1.29560e-03'
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_0 = '3.09406e-03*lvn_subvt*lvn_subvt+-1.23763e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_1 = '3.10416e-03*lvn_subvt*lvn_subvt+1.24166e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0 = '1.10588e+03*lvn_saturation*lvn_saturation+9.76162e+03*lvn_saturation+3.85540e+03'
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1 = '-6.14031e+02*lvn_saturation*lvn_saturation+3.55288e+03*lvn_saturation+1.36790e+04'
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0 = '-2.37156e-04*lvn_threshold*lvn_threshold+5.41889e-02*lvn_threshold+-1.56630e-01'
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1 = '-3.54442e-03*lvn_threshold*lvn_threshold+4.54875e-02*lvn_threshold+-5.70930e-03'
+ sky130_fd_pr__special_nfet_pass_flash__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult = '2.36250e-04*hvtox*hvtox+3.48425e-02*hvtox+8.98050e-01'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult = '1.87500e-06*hvn_diode*hvn_diode+5.91425e-02*hvn_diode+1.01440e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult = '5.00000e-02*hvn_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0 = '6.73731e-05*hvn_bodyeffect*hvn_bodyeffect+1.44721e-03*hvn_bodyeffect+5.94980e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1 = '4.82875e-05*hvn_bodyeffect*hvn_bodyeffect+2.60342e-03*hvn_bodyeffect+-6.80590e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2 = '5.88812e-05*hvn_bodyeffect*hvn_bodyeffect+1.91960e-03*hvn_bodyeffect+-1.71730e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0 = '-7.68594e-05*hvn_mobility*hvn_mobility+1.74013e-04*hvn_mobility+-1.64490e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1 = '-6.29875e-05*hvn_mobility*hvn_mobility+3.40150e-04*hvn_mobility+-2.93900e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2 = '-1.05841e-04*hvn_mobility*hvn_mobility+-8.23638e-04*hvn_mobility+-4.10540e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0 = '-1.58063e+01*hvn_saturation*hvn_saturation+2.77575e+03*hvn_saturation+1.10090e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1 = '-1.25478e+02*hvn_saturation*hvn_saturation+1.14561e+03*hvn_saturation+-3.86290e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2 = '1.89456e+02*hvn_saturation*hvn_saturation+3.27588e+03*hvn_saturation+-5.55680e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0 = '-1.66438e-04*hvn_threshold*hvn_threshold+1.97085e-02*hvn_threshold+-1.50750e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1 = '-1.62219e-04*hvn_threshold*hvn_threshold+1.69419e-02*hvn_threshold+-1.26710e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2 = '-1.69625e-04*hvn_threshold*hvn_threshold+1.76940e-02*hvn_threshold+-2.21230e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0 = '6.49969e-05*hvn_bodyeffect*hvn_bodyeffect+1.48076e-03*hvn_bodyeffect+1.31270e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1 = '4.33569e-05*hvn_bodyeffect*hvn_bodyeffect+2.97512e-03*hvn_bodyeffect+-5.34210e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0 = '-7.58844e-05*hvn_mobility*hvn_mobility+2.36187e-04*hvn_mobility+-2.96850e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1 = '-5.67477e-05*hvn_mobility*hvn_mobility+5.00359e-04*hvn_mobility+-1.01150e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0 = '-1.05934e+02*hvn_saturation*hvn_saturation+1.86891e+03*hvn_saturation+-3.50340e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1 = '-1.37866e+02*hvn_saturation*hvn_saturation+1.07262e+03*hvn_saturation+3.23350e+02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0 = '-1.63406e-04*hvn_threshold*hvn_threshold+1.97464e-02*hvn_threshold+-1.52620e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1 = '-1.63219e-04*hvn_threshold*hvn_threshold+1.69772e-02*hvn_threshold+-2.53650e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0 = '6.42844e-05*hvn_bodyeffect*hvn_bodyeffect+1.50469e-03*hvn_bodyeffect+1.01730e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1 = '4.41862e-05*hvn_bodyeffect*hvn_bodyeffect+2.84487e-03*hvn_bodyeffect+-5.78480e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2 = '5.32719e-05*hvn_bodyeffect*hvn_bodyeffect+2.20489e-03*hvn_bodyeffect+-1.51370e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0 = '-7.63000e-05*hvn_mobility*hvn_mobility+2.03675e-04*hvn_mobility+-3.12710e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1 = '-5.58209e-05*hvn_mobility*hvn_mobility+4.70666e-04*hvn_mobility+-1.39930e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2 = '-6.19250e-05*hvn_mobility*hvn_mobility+3.00125e-04*hvn_mobility+-3.00200e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0 = '-8.86719e+01*hvn_saturation*hvn_saturation+1.90121e+03*hvn_saturation+-3.94640e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1 = '-1.36300e+02*hvn_saturation*hvn_saturation+1.00510e+03*hvn_saturation+-1.84170e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2 = '-1.28133e+02*hvn_saturation*hvn_saturation+1.10697e+03*hvn_saturation+-2.99490e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0 = '-1.63094e-04*hvn_threshold*hvn_threshold+1.96286e-02*hvn_threshold+-2.45260e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1 = '-1.60731e-04*hvn_threshold*hvn_threshold+1.69806e-02*hvn_threshold+-9.99980e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2 = '-1.61125e-04*hvn_threshold*hvn_threshold+1.79651e-02*hvn_threshold+-8.21650e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult = '3.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42 = '3.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult = '3.12500e-03*nfet_01v8_lvt*nfet_01v8_lvt+7.50000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42 = '8.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult = '3.12500e-03*lvln_mobility*lvln_mobility+7.50000e-02*lvln_mobility+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42 = '8.75000e-02*lvln_mobility+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult = '-2.59375e-05*lvn_diode*lvn_diode+4.38787e-02*lvn_diode+1.00040e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff = '-4.91625e-11*poly_cd*poly_cd+-3.37112e-09*poly_cd+-1.36190e-09'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult = '-2.39062e-04*lvtox*lvtox+1.49487e-02*lvtox+9.24290e-01'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult = '4.43125e-04*lvn_diode*lvn_diode+3.72125e-02*lvn_diode+8.91760e-01'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult = '5.00000e-02*lvln_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0 = '2.16537e-04*lvln_bodyeffect*lvln_bodyeffect+-2.62240e-03*lvln_bodyeffect+-1.78380e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1 = '1.35078e-04*lvln_bodyeffect*lvln_bodyeffect+-2.77109e-03*lvln_bodyeffect+-8.88490e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2 = '2.44556e-05*lvln_bodyeffect*lvln_bodyeffect+4.77047e-04*lvln_bodyeffect+-1.89470e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3 = '3.99562e-04*lvln_bodyeffect*lvln_bodyeffect+-5.82675e-03*lvln_bodyeffect+-1.30740e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4 = '1.72656e-04*lvln_bodyeffect*lvln_bodyeffect+-4.12787e-03*lvln_bodyeffect+-8.65900e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5 = '5.23656e-05*lvln_bodyeffect*lvln_bodyeffect+-1.42609e-03*lvln_bodyeffect+-1.49170e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6 = '2.87944e-04*lvln_bodyeffect*lvln_bodyeffect+-4.77777e-03*lvln_bodyeffect+-2.04570e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7 = '1.70841e-04*lvln_bodyeffect*lvln_bodyeffect+-3.84876e-03*lvln_bodyeffect+-9.14240e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8 = '4.93312e-05*lvln_bodyeffect*lvln_bodyeffect+-1.29807e-03*lvln_bodyeffect+-1.35180e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0 = '-1.27475e-05*lvln_mobility*lvln_mobility+-3.77012e-04*lvln_mobility+-2.59890e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1 = '-3.12666e-05*lvln_mobility*lvln_mobility+-1.65496e-04*lvln_mobility+6.88700e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2 = '-3.05450e-05*lvln_mobility*lvln_mobility+-3.54088e-04*lvln_mobility+7.01070e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3 = '-2.20438e-05*lvln_mobility*lvln_mobility+-1.72850e-04*lvln_mobility+-4.13870e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4 = '-2.53094e-05*lvln_mobility*lvln_mobility+2.66612e-04*lvln_mobility+-2.15790e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5 = '-2.68078e-05*lvln_mobility*lvln_mobility+-3.03044e-04*lvln_mobility+-1.04250e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6 = '-2.88062e-05*lvln_mobility*lvln_mobility+1.33150e-04*lvln_mobility+-8.36300e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7 = '-2.50531e-05*lvln_mobility*lvln_mobility+1.44313e-04*lvln_mobility+-4.23970e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8 = '-2.64838e-05*lvln_mobility*lvln_mobility+-4.36215e-04*lvln_mobility+-1.91930e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0 = '7.32625e+01*lvln_saturation*lvln_saturation+7.38425e+03*lvln_saturation+-4.14020e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1 = '2.23044e+02*lvln_saturation*lvln_saturation+7.08838e+03*lvln_saturation+-1.70920e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2 = '1.66750e+02*lvln_saturation*lvln_saturation+4.82325e+03*lvln_saturation+-3.89100e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3 = '1.01919e+02*lvln_saturation*lvln_saturation+8.30375e+03*lvln_saturation+-6.08870e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4 = '7.99125e+01*lvln_saturation*lvln_saturation+6.43850e+03*lvln_saturation+-1.51960e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5 = '2.15024e+02*lvln_saturation*lvln_saturation+5.42662e+03*lvln_saturation+-4.15880e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6 = '-5.46875e+00*lvln_saturation*lvln_saturation+6.40075e+03*lvln_saturation+-5.55550e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7 = '8.60469e+01*lvln_saturation*lvln_saturation+5.73812e+03*lvln_saturation+-7.90250e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8 = '3.04746e+02*lvln_saturation*lvln_saturation+5.30988e+03*lvln_saturation+-1.05440e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0 = '-2.61075e-04*lvln_threshold*lvln_threshold+1.48638e-02*lvln_threshold+-1.90980e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1 = '-1.89812e-04*lvln_threshold*lvln_threshold+1.33500e-02*lvln_threshold+-2.59700e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2 = '-8.61250e-05*lvln_threshold*lvln_threshold+7.26675e-03*lvln_threshold+-1.23440e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3 = '-4.21469e-04*lvln_threshold*lvln_threshold+1.39709e-02*lvln_threshold+-1.12620e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4 = '-2.22750e-04*lvln_threshold*lvln_threshold+1.09125e-02*lvln_threshold+-2.00030e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5 = '-9.39187e-05*lvln_threshold*lvln_threshold+5.23312e-03*lvln_threshold+-7.42980e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6 = '-3.57906e-04*lvln_threshold*lvln_threshold+1.21069e-02*lvln_threshold+-1.02570e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7 = '-2.25563e-04*lvln_threshold*lvln_threshold+9.05225e-03*lvln_threshold+-1.70600e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8 = '-9.28219e-05*lvln_threshold*lvln_threshold+4.10981e-03*lvln_threshold+-6.94560e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0 = '2.12059e-04*lvln_bodyeffect*lvln_bodyeffect+-2.43399e-03*lvln_bodyeffect+-1.75260e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1 = '1.29553e-04*lvln_bodyeffect*lvln_bodyeffect+-2.65451e-03*lvln_bodyeffect+-9.39780e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2 = '4.61625e-05*lvln_bodyeffect*lvln_bodyeffect+-1.24362e-03*lvln_bodyeffect+-2.33740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3 = '3.91781e-04*lvln_bodyeffect*lvln_bodyeffect+-5.71988e-03*lvln_bodyeffect+-1.42820e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4 = '1.47672e-04*lvln_bodyeffect*lvln_bodyeffect+-3.83104e-03*lvln_bodyeffect+-9.64160e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5 = '4.74750e-05*lvln_bodyeffect*lvln_bodyeffect+-1.34908e-03*lvln_bodyeffect+-2.71180e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6 = '3.32397e-04*lvln_bodyeffect*lvln_bodyeffect+-5.34884e-03*lvln_bodyeffect+-1.91600e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7 = '1.37456e-04*lvln_bodyeffect*lvln_bodyeffect+-3.47033e-03*lvln_bodyeffect+-1.14380e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8 = '4.66500e-05*lvln_bodyeffect*lvln_bodyeffect+-1.20602e-03*lvln_bodyeffect+-2.83740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0 = '-1.76219e-05*lvln_mobility*lvln_mobility+-2.84613e-04*lvln_mobility+-6.03480e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1 = '-3.21063e-05*lvln_mobility*lvln_mobility+-6.38750e-05*lvln_mobility+-2.81360e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2 = '-2.79550e-05*lvln_mobility*lvln_mobility+-3.72130e-04*lvln_mobility+-1.72530e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3 = '-2.89937e-05*lvln_mobility*lvln_mobility+-9.04500e-05*lvln_mobility+-4.67570e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4 = '-2.23969e-05*lvln_mobility*lvln_mobility+2.08213e-04*lvln_mobility+-6.94280e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5 = '-2.35313e-05*lvln_mobility*lvln_mobility+-2.96250e-04*lvln_mobility+-4.24740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6 = '-3.00687e-05*lvln_mobility*lvln_mobility+1.03425e-04*lvln_mobility+-6.15790e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7 = '-2.47250e-05*lvln_mobility*lvln_mobility+5.17000e-05*lvln_mobility+-8.45140e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8 = '-2.26906e-05*lvln_mobility*lvln_mobility+-4.28638e-04*lvln_mobility+-6.56350e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0 = '1.74569e+02*lvln_saturation*lvln_saturation+7.96162e+03*lvln_saturation+1.45400e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1 = '2.40744e+02*lvln_saturation*lvln_saturation+7.13262e+03*lvln_saturation+-1.62240e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2 = '1.56794e+02*lvln_saturation*lvln_saturation+5.01475e+03*lvln_saturation+2.32830e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3 = '1.09244e+02*lvln_saturation*lvln_saturation+8.25900e+03*lvln_saturation+-6.71990e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4 = '1.60491e+02*lvln_saturation*lvln_saturation+6.83362e+03*lvln_saturation+3.27640e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5 = '3.10119e+02*lvln_saturation*lvln_saturation+5.98098e+03*lvln_saturation+9.08320e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6 = '6.03562e+01*lvln_saturation*lvln_saturation+7.56138e+03*lvln_saturation+-6.43120e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7 = '1.54125e+02*lvln_saturation*lvln_saturation+6.14912e+03*lvln_saturation+-2.62550e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8 = '5.30047e+02*lvln_saturation*lvln_saturation+7.52931e+03*lvln_saturation+1.41900e+04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0 = '-2.69669e-04*lvln_threshold*lvln_threshold+1.48915e-02*lvln_threshold+-5.11330e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1 = '-1.94688e-04*lvln_threshold*lvln_threshold+1.34505e-02*lvln_threshold+-1.00420e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2 = '-8.10625e-05*lvln_threshold*lvln_threshold+7.25900e-03*lvln_threshold+-1.77560e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3 = '-4.34213e-04*lvln_threshold*lvln_threshold+1.42046e-02*lvln_threshold+-8.51510e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4 = '-1.97313e-04*lvln_threshold*lvln_threshold+1.04557e-02*lvln_threshold+-1.70880e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5 = '-8.34781e-05*lvln_threshold*lvln_threshold+4.97284e-03*lvln_threshold+-1.99910e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6 = '-3.76781e-04*lvln_threshold*lvln_threshold+1.26681e-02*lvln_threshold+-1.30210e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7 = '-1.85438e-04*lvln_threshold*lvln_threshold+8.48675e-03*lvln_threshold+-1.86740e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8 = '-8.59000e-05*lvln_threshold*lvln_threshold+3.90465e-03*lvln_threshold+-2.40190e-02'
+ sky130_fd_pr__special_nfet_pass_lvt__ajunction_mult = '-2.59375e-05*lvn_diode*lvn_diode+4.38787e-02*lvn_diode+1.00040e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__dlc_diff = '-4.91625e-11*poly_cd*poly_cd+3.37112e-09*poly_cd+-1.36190e-09'
+ sky130_fd_pr__special_nfet_pass_lvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass_lvt__lint_diff = '4.33125e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_lvt__nfactor_diff_0 = '-2.46134e-02*lvn_subvt*lvn_subvt+1.00321e-01*lvn_subvt+3.97550e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__overlap_mult = '-2.39062e-04*lvtox*lvtox+1.49487e-02*lvtox+9.24290e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult = '4.43125e-04*lvn_diode*lvn_diode+3.72125e-02*lvn_diode+8.91760e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__rshn_mult = '5.00000e-02*special_nfet_pass_lvt+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__u0_diff_0 = '-3.63906e-05*lvln_mobility*lvln_mobility+3.15216e-03*lvln_mobility+-6.97310e-03'
+ sky130_fd_pr__special_nfet_pass_lvt__vsat_diff_0 = '6.84562e+01*lvln_saturation*lvln_saturation+1.18361e+04*lvln_saturation+8.11120e+03'
+ sky130_fd_pr__special_nfet_pass_lvt__vth0_diff_0 = '5.66969e-04*lvln_threshold*lvln_threshold+3.27404e-02*lvln_threshold+2.47670e-02'
+ sky130_fd_pr__special_nfet_pass_lvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_pass__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass__overlap_mult = '-1.27188e-04*lvtox*lvtox+8.00875e-03*lvtox+9.84200e-01'
+ sky130_fd_pr__special_nfet_pass__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_pass__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass__u0_diff_0 = '3.55678e-04*lvn_mobility*lvn_mobility+3.05794e-03*lvn_mobility+-2.92260e-03'
+ sky130_fd_pr__special_nfet_pass__vth0_diff_0 = '-2.68250e-04*lvn_threshold*lvn_threshold+4.27650e-02*lvn_threshold+2.75220e-02'
+ sky130_fd_pr__special_nfet_pass__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_latch__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_latch__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_latch__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_latch__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_latch__overlap_mult = '-1.27188e-04*lvtox*lvtox+8.00875e-03*lvtox+9.84200e-01'
+ sky130_fd_pr__special_nfet_latch__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_latch__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_latch__u0_diff_0 = '6.25750e-06*lvn_mobility*lvn_mobility+2.32240e-03*lvn_mobility+3.03680e-04'
+ sky130_fd_pr__special_nfet_latch__vth0_diff_0 = '-9.35625e-05*lvn_threshold*lvn_threshold+3.22038e-02*lvn_threshold+2.09520e-02'
+ sky130_fd_pr__special_nfet_latch__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult = '-1.87500e-06*lvn_diode*lvn_diode+5.53750e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__rf_nfet_01v8_b__dlc_diff = '-1.06849e-10*poly_cd*poly_cd+-3.77438e-09*poly_cd+-6.14920e-10'
+ sky130_fd_pr__rf_nfet_01v8_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_01v8_b__overlap_mult = '-6.32500e-04*lvtox*lvtox+1.48000e-03*lvtox+9.64200e-01'
+ sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult = '-1.25000e-06*lvn_diode*lvn_diode+5.67550e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult = '5.00000e-02*lvn_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_01v8_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_0 = '9.86813e-05*lvn_bodyeffect*lvn_bodyeffect+-2.16475e-04*lvn_bodyeffect+7.64020e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_1 = '3.98437e-05*lvn_bodyeffect*lvn_bodyeffect+-8.01375e-04*lvn_bodyeffect+1.68400e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_2 = '2.04688e-05*lvn_bodyeffect*lvn_bodyeffect+-7.86125e-04*lvn_bodyeffect+3.45610e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_3 = '1.15172e-04*lvn_bodyeffect*lvn_bodyeffect+-1.04921e-03*lvn_bodyeffect+4.58640e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_4 = '8.01562e-05*lvn_bodyeffect*lvn_bodyeffect+-2.15937e-03*lvn_bodyeffect+2.04550e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_5 = '3.81250e-05*lvn_bodyeffect*lvn_bodyeffect+-1.28100e-03*lvn_bodyeffect+3.72450e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_6 = '1.12641e-04*lvn_bodyeffect*lvn_bodyeffect+-6.86062e-04*lvn_bodyeffect+1.94870e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_7 = '7.50000e-05*lvn_bodyeffect*lvn_bodyeffect+-1.86975e-03*lvn_bodyeffect+1.77710e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_8 = '3.85937e-05*lvn_bodyeffect*lvn_bodyeffect+-1.41812e-03*lvn_bodyeffect+3.54600e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_0 = '-2.03169e-05*lvn_mobility*lvn_mobility+-7.14350e-05*lvn_mobility+7.86820e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_1 = '-2.40125e-05*lvn_mobility*lvn_mobility+-2.04582e-04*lvn_mobility+6.95070e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_2 = '-2.55544e-05*lvn_mobility*lvn_mobility+-3.10587e-04*lvn_mobility+-1.86680e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_3 = '-1.55000e-05*lvn_mobility*lvn_mobility+-4.14350e-04*lvn_mobility+-5.08880e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_4 = '-2.01469e-05*lvn_mobility*lvn_mobility+-9.54875e-05*lvn_mobility+-3.38250e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_5 = '-2.12863e-05*lvn_mobility*lvn_mobility+-3.87613e-04*lvn_mobility+-1.08370e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_6 = '-1.66125e-05*lvn_mobility*lvn_mobility+-1.83325e-04*lvn_mobility+-3.81310e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_7 = '-1.86562e-05*lvn_mobility*lvn_mobility+-7.10500e-05*lvn_mobility+-3.65260e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_8 = '-2.01562e-05*lvn_mobility*lvn_mobility+-3.97775e-04*lvn_mobility+-2.32590e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_0 = '-1.15489e+02*lvn_saturation*lvn_saturation+5.36138e+03*lvn_saturation+8.76330e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_1 = '4.23912e+01*lvn_saturation*lvn_saturation+5.05100e+03*lvn_saturation+2.92740e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_2 = '2.37344e+02*lvn_saturation*lvn_saturation+6.14662e+03*lvn_saturation+4.00800e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_3 = '-1.44812e+01*lvn_saturation*lvn_saturation+5.13850e+03*lvn_saturation+-7.67730e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_4 = '1.45662e+02*lvn_saturation*lvn_saturation+6.06888e+03*lvn_saturation+-3.22610e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_5 = '2.18925e+02*lvn_saturation*lvn_saturation+5.16400e+03*lvn_saturation+-3.10380e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_6 = '-1.10087e+02*lvn_saturation*lvn_saturation+4.09440e+03*lvn_saturation+-1.05210e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_7 = '1.07662e+02*lvn_saturation*lvn_saturation+5.22625e+03*lvn_saturation+-3.85660e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_8 = '1.96437e+02*lvn_saturation*lvn_saturation+4.60912e+03*lvn_saturation+-7.49490e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_0 = '-1.62094e-04*lvn_threshold*lvn_threshold+1.35881e-02*lvn_threshold+-1.90450e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_1 = '-7.34188e-05*lvn_threshold*lvn_threshold+8.96013e-03*lvn_threshold+-2.47180e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_2 = '-4.36562e-05*lvn_threshold*lvn_threshold+7.71487e-03*lvn_threshold+-1.14640e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_3 = '-1.64381e-04*lvn_threshold*lvn_threshold+8.90112e-03*lvn_threshold+3.12960e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_4 = '-1.15569e-04*lvn_threshold*lvn_threshold+7.71322e-03*lvn_threshold+-1.91180e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_5 = '-5.94469e-05*lvn_threshold*lvn_threshold+5.11071e-03*lvn_threshold+-1.09280e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_6 = '-1.75688e-04*lvn_threshold*lvn_threshold+7.06775e-03*lvn_threshold+-1.03570e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_7 = '-1.04675e-04*lvn_threshold*lvn_threshold+6.36330e-03*lvn_threshold+-1.86330e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_8 = '-5.97938e-05*lvn_threshold*lvn_threshold+4.31957e-03*lvn_threshold+-1.47380e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_0 = '1.01206e-04*lvn_bodyeffect*lvn_bodyeffect+-2.39325e-04*lvn_bodyeffect+6.60760e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_1 = '7.19375e-05*lvn_bodyeffect*lvn_bodyeffect+-1.34700e-03*lvn_bodyeffect+2.24380e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_2 = '3.36875e-05*lvn_bodyeffect*lvn_bodyeffect+-1.03250e-03*lvn_bodyeffect+3.75000e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_3 = '1.50000e-04*lvn_bodyeffect*lvn_bodyeffect+-1.47690e-03*lvn_bodyeffect+5.54840e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_4 = '9.85312e-05*lvn_bodyeffect*lvn_bodyeffect+-2.44437e-03*lvn_bodyeffect+2.36230e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_5 = '4.27812e-05*lvn_bodyeffect*lvn_bodyeffect+-1.40612e-03*lvn_bodyeffect+3.90920e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_6 = '1.46059e-04*lvn_bodyeffect*lvn_bodyeffect+-1.06724e-03*lvn_bodyeffect+2.99510e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_7 = '9.85000e-05*lvn_bodyeffect*lvn_bodyeffect+-2.19400e-03*lvn_bodyeffect+2.15790e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_8 = '4.26875e-05*lvn_bodyeffect*lvn_bodyeffect+-1.52550e-03*lvn_bodyeffect+3.73290e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_0 = '-2.36125e-05*lvn_mobility*lvn_mobility+-9.13050e-05*lvn_mobility+-6.96680e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_1 = '-2.69156e-05*lvn_mobility*lvn_mobility+-1.03337e-04*lvn_mobility+-1.34750e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_2 = '-2.58159e-05*lvn_mobility*lvn_mobility+-2.66011e-04*lvn_mobility+-1.00130e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_3 = '-1.96437e-05*lvn_mobility*lvn_mobility+-3.09800e-04*lvn_mobility+-5.73800e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_4 = '-2.20062e-05*lvn_mobility*lvn_mobility+1.62250e-05*lvn_mobility+-6.72530e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_5 = '-2.11250e-05*lvn_mobility*lvn_mobility+-2.42950e-04*lvn_mobility+-4.97740e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_6 = '-1.91562e-05*lvn_mobility*lvn_mobility+-1.70875e-04*lvn_mobility+-3.71750e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_7 = '-2.06969e-05*lvn_mobility*lvn_mobility+4.18625e-05*lvn_mobility+-5.53610e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_8 = '-2.02562e-05*lvn_mobility*lvn_mobility+-3.29650e-04*lvn_mobility+-4.09270e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_0 = '-6.86938e+01*lvn_saturation*lvn_saturation+5.32662e+03*lvn_saturation+-9.57840e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_1 = '1.42819e+02*lvn_saturation*lvn_saturation+5.97550e+03*lvn_saturation+-1.94710e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_2 = '4.07231e+02*lvn_saturation*lvn_saturation+7.37000e+03*lvn_saturation+3.93430e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_3 = '-1.55125e+01*lvn_saturation*lvn_saturation+5.34838e+03*lvn_saturation+-9.28630e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_4 = '2.14356e+02*lvn_saturation*lvn_saturation+6.49375e+03*lvn_saturation+-2.37570e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_5 = '5.62681e+02*lvn_saturation*lvn_saturation+7.95552e+03*lvn_saturation+1.42910e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_6 = '-1.00753e+02*lvn_saturation*lvn_saturation+4.25624e+03*lvn_saturation+-1.13210e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_7 = '7.49312e+01*lvn_saturation*lvn_saturation+4.89662e+03*lvn_saturation+-8.60840e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_8 = '5.51006e+02*lvn_saturation*lvn_saturation+7.46000e+03*lvn_saturation+9.12790e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_0 = '-1.63794e-04*lvn_threshold*lvn_threshold+1.35991e-02*lvn_threshold+5.51620e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_1 = '-1.14875e-04*lvn_threshold*lvn_threshold+9.79050e-03*lvn_threshold+-1.71250e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_2 = '-6.13437e-05*lvn_threshold*lvn_threshold+8.03163e-03*lvn_threshold+-1.35250e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_3 = '-2.02750e-04*lvn_threshold*lvn_threshold+9.64162e-03*lvn_threshold+-5.00650e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_4 = '-1.44725e-04*lvn_threshold*lvn_threshold+8.33085e-03*lvn_threshold+-2.55090e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_5 = '-6.63719e-05*lvn_threshold*lvn_threshold+5.42226e-03*lvn_threshold+-1.84290e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_6 = '-2.01062e-04*lvn_threshold*lvn_threshold+7.62525e-03*lvn_threshold+-1.13020e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_7 = '-1.45200e-04*lvn_threshold*lvn_threshold+7.05445e-03*lvn_threshold+-2.98950e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_8 = '-6.84031e-05*lvn_threshold*lvn_threshold+4.64789e-03*lvn_threshold+-1.92140e-02'
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult = '3.75000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2 = '3.75000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult = '6.87500e-03*pfet_01v8*pfet_01v8+8.50000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2 = '3.12500e-03*pfet_01v8*pfet_01v8+6.25000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult = '6.87500e-03*lvp_mobility*lvp_mobility+8.50000e-02*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2 = '3.12500e-03*lvp_mobility*lvp_mobility+6.25000e-02*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult = '-3.12500e-07*lvp_diode*lvp_diode+2.36612e-02*lvp_diode+9.96260e-01'
+ sky130_fd_pr__rf_pfet_01v8_b__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__overlap_mult = '7.47062e-03*lvtox*lvtox+2.98800e-02*lvtox+9.54350e-01'
+ sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult = '2.18750e-06*lvp_diode*lvp_diode+2.37662e-02*lvp_diode+1.00090e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult = '5.00000e-02*lvp_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_pfet_01v8_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0 = '7.88925e-04*lvp_bodyeffect*lvp_bodyeffect+-3.74695e-03*lvp_bodyeffect+-2.39530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1 = '4.12838e-04*lvp_bodyeffect*lvp_bodyeffect+-7.85000e-05*lvp_bodyeffect+-1.46000e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2 = '8.07491e-05*lvp_bodyeffect*lvp_bodyeffect+4.28325e-03*lvp_bodyeffect+-1.75040e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3 = '8.30297e-04*lvp_bodyeffect*lvp_bodyeffect+-2.77369e-03*lvp_bodyeffect+-2.56720e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4 = '4.43511e-04*lvp_bodyeffect*lvp_bodyeffect+-2.39504e-03*lvp_bodyeffect+-1.64290e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5 = '1.27375e-04*lvp_bodyeffect*lvp_bodyeffect+1.05000e-05*lvp_bodyeffect+-1.85780e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6 = '8.48497e-04*lvp_bodyeffect*lvp_bodyeffect+-2.83474e-03*lvp_bodyeffect+-2.63870e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7 = '4.38997e-04*lvp_bodyeffect*lvp_bodyeffect+-1.75149e-03*lvp_bodyeffect+-1.36950e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8 = '1.16562e-04*lvp_bodyeffect*lvp_bodyeffect+8.99500e-04*lvp_bodyeffect+-1.78310e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0 = '-2.95281e-06*lvp_mobility*lvp_mobility+1.07038e-05*lvp_mobility+-2.56080e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1 = '-3.17469e-06*lvp_mobility*lvp_mobility+-7.32625e-06*lvp_mobility+-1.75340e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2 = '-5.07816e-06*lvp_mobility*lvp_mobility+-4.14349e-05*lvp_mobility+-1.15280e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3 = '-1.61219e-06*lvp_mobility*lvp_mobility+-4.63037e-05*lvp_mobility+-4.39530e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4 = '-2.81625e-06*lvp_mobility*lvp_mobility+-8.32000e-06*lvp_mobility+-4.02980e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5 = '-3.43469e-06*lvp_mobility*lvp_mobility+-2.94162e-05*lvp_mobility+-2.29660e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6 = '-1.04187e-06*lvp_mobility*lvp_mobility+-6.76675e-05*lvp_mobility+-7.89060e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7 = '-3.19031e-06*lvp_mobility*lvp_mobility+-2.56063e-05*lvp_mobility+-3.06110e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8 = '-2.76312e-06*lvp_mobility*lvp_mobility+-4.04825e-05*lvp_mobility+-3.26940e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0 = '-2.19959e+02*lvp_saturation*lvp_saturation+3.58099e+03*lvp_saturation+-1.79270e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1 = '-6.67469e+02*lvp_saturation*lvp_saturation+2.31875e+02*lvp_saturation+-3.93900e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2 = '-3.74053e+02*lvp_saturation*lvp_saturation+-8.13988e+02*lvp_saturation+-3.70520e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3 = '-4.49481e+02*lvp_saturation*lvp_saturation+9.72500e+02*lvp_saturation+-7.60430e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4 = '-5.17684e+02*lvp_saturation*lvp_saturation+8.18238e+02*lvp_saturation+2.22900e+02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5 = '-1.04765e+03*lvp_saturation*lvp_saturation+-8.24300e+02*lvp_saturation+1.23580e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6 = '-5.68250e+02*lvp_saturation*lvp_saturation+8.48900e+02*lvp_saturation+-3.99640e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7 = '-6.26394e+02*lvp_saturation*lvp_saturation+6.40750e+02*lvp_saturation+-5.40770e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8 = '-8.45866e+02*lvp_saturation*lvp_saturation+-1.39554e+03*lvp_saturation+2.23200e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0 = '-2.08957e-03*lvp_threshold*lvp_threshold+1.60973e-02*lvp_threshold+5.41510e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1 = '-1.03035e-03*lvp_threshold*lvp_threshold+1.53896e-02*lvp_threshold+-1.32890e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2 = '-2.39119e-04*lvp_threshold*lvp_threshold+6.98988e-03*lvp_threshold+1.68740e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3 = '-2.17209e-03*lvp_threshold*lvp_threshold+2.30241e-02*lvp_threshold+5.54000e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4 = '-1.09537e-03*lvp_threshold*lvp_threshold+1.57754e-02*lvp_threshold+9.01640e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5 = '-2.77719e-04*lvp_threshold*lvp_threshold+6.42650e-03*lvp_threshold+4.31850e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6 = '-2.17009e-03*lvp_threshold*lvp_threshold+2.74224e-02*lvp_threshold+1.32910e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7 = '-1.05824e-03*lvp_threshold*lvp_threshold+1.65510e-02*lvp_threshold+5.46190e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8 = '-2.81481e-04*lvp_threshold*lvp_threshold+8.40712e-03*lvp_threshold+3.05520e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0 = '8.11859e-04*lvp_bodyeffect*lvp_bodyeffect+-3.96794e-03*lvp_bodyeffect+-2.22710e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1 = '4.22813e-04*lvp_bodyeffect*lvp_bodyeffect+-2.25700e-04*lvp_bodyeffect+-1.40490e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2 = '7.11859e-05*lvp_bodyeffect*lvp_bodyeffect+4.23974e-03*lvp_bodyeffect+-1.85950e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3 = '8.25749e-04*lvp_bodyeffect*lvp_bodyeffect+-2.75950e-03*lvp_bodyeffect+-2.34610e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4 = '4.42350e-04*lvp_bodyeffect*lvp_bodyeffect+-2.42190e-03*lvp_bodyeffect+-1.27890e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5 = '1.26969e-04*lvp_bodyeffect*lvp_bodyeffect+-2.36250e-05*lvp_bodyeffect+-1.85990e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6 = '8.47931e-04*lvp_bodyeffect*lvp_bodyeffect+-2.95897e-03*lvp_bodyeffect+-2.51000e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7 = '4.38387e-04*lvp_bodyeffect*lvp_bodyeffect+-1.69255e-03*lvp_bodyeffect+-1.09530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8 = '1.15937e-04*lvp_bodyeffect*lvp_bodyeffect+8.62750e-04*lvp_bodyeffect+-1.66060e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0 = '-3.02500e-06*lvp_mobility*lvp_mobility+6.14500e-06*lvp_mobility+-4.34040e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1 = '-3.78563e-06*lvp_mobility*lvp_mobility+-1.01825e-05*lvp_mobility+-2.53300e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2 = '-3.14672e-06*lvp_mobility*lvp_mobility+-4.08281e-05*lvp_mobility+-1.85700e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3 = '-5.81562e-07*lvp_mobility*lvp_mobility+-4.06338e-05*lvp_mobility+-5.35030e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4 = '-2.25750e-06*lvp_mobility*lvp_mobility+-1.96525e-05*lvp_mobility+-6.24650e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5 = '-3.40312e-06*lvp_mobility*lvp_mobility+-3.32025e-05*lvp_mobility+-3.34450e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6 = '-7.05625e-07*lvp_mobility*lvp_mobility+-7.59700e-05*lvp_mobility+-6.46020e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7 = '-3.02000e-06*lvp_mobility*lvp_mobility+-2.82000e-05*lvp_mobility+-5.75480e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8 = '-2.91781e-06*lvp_mobility*lvp_mobility+-4.52087e-05*lvp_mobility+-4.40410e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0 = '-3.93106e+02*lvp_saturation*lvp_saturation+3.06255e+03*lvp_saturation+-1.65610e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1 = '-4.90413e+02*lvp_saturation*lvp_saturation+1.33069e+03*lvp_saturation+8.76350e+02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2 = '-1.32498e+03*lvp_saturation*lvp_saturation+-1.38783e+03*lvp_saturation+1.59210e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3 = '-6.36825e+02*lvp_saturation*lvp_saturation+7.42250e+02*lvp_saturation+-2.98080e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4 = '-6.15031e+02*lvp_saturation*lvp_saturation+1.22375e+02*lvp_saturation+-1.15500e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5 = '-1.24004e+03*lvp_saturation*lvp_saturation+-8.54950e+02*lvp_saturation+9.11750e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6 = '-5.66359e+02*lvp_saturation*lvp_saturation+1.15776e+03*lvp_saturation+-2.85020e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7 = '-6.28938e+02*lvp_saturation*lvp_saturation+3.11750e+02*lvp_saturation+-3.91400e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8 = '-1.01133e+03*lvp_saturation*lvp_saturation+-2.22694e+03*lvp_saturation+1.14100e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0 = '-2.10059e-03*lvp_threshold*lvp_threshold+1.63614e-02*lvp_threshold+1.80470e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1 = '-1.01603e-03*lvp_threshold*lvp_threshold+1.54661e-02*lvp_threshold+1.24260e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2 = '-2.85394e-04*lvp_threshold*lvp_threshold+6.92225e-03*lvp_threshold+9.47730e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3 = '-2.19548e-03*lvp_threshold*lvp_threshold+2.26099e-02*lvp_threshold+6.48720e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4 = '-1.11394e-03*lvp_threshold*lvp_threshold+1.57338e-02*lvp_threshold+2.23420e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5 = '-2.83188e-04*lvp_threshold*lvp_threshold+6.39900e-03*lvp_threshold+1.20970e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6 = '-2.17306e-03*lvp_threshold*lvp_threshold+2.71660e-02*lvp_threshold+1.77530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7 = '-1.05896e-03*lvp_threshold*lvp_threshold+1.65740e-02*lvp_threshold+9.71640e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8 = '-2.80031e-04*lvp_threshold*lvp_threshold+8.37688e-03*lvp_threshold+1.54910e-02'
+ rcl1 = '1.75000e-01*ic_res*ic_res+2.62500e+00*ic_res+9.30000e+00'
+ rcn = '1.59375e+00*ic_res_ndiff*ic_res_ndiff+3.43750e+01*ic_res_ndiff+1.82000e+02'
+ rcp = '6.75000e+01*ic_res_pdiff+6.00000e+02'
+ rcp1 = '-6.87500e-01*ic_res_poly*ic_res_poly+2.72500e+01*ic_res_poly+1.45280e+02'
+ rcvia = '2.50000e-01*ic_res*ic_res+1.62500e+00*ic_res+4.50000e+00'
+ rcvia2 = '5.25000e-02*ic_res*ic_res+9.37500e-01*ic_res+3.41000e+00'
+ rcvia3 = '5.25000e-02*ic_res*ic_res+9.37500e-01*ic_res+3.41000e+00'
+ rcvia4 = '4.46875e-03*ic_res*ic_res+1.09875e-01*ic_res+3.80000e-01'
+ rdn_hv = '3.00000e+00*ic_res_ndiff+1.14000e+02'
+ rdp_hv = '7.75000e+00*ic_res_pdiff+1.91000e+02'
+ rl1 = '-3.12500e-03*ic_res*ic_res+6.62500e-01*ic_res+1.22000e+01'
+ rm1 = '5.00000e-03*ic_res+1.25000e-01'
+ rm2 = '5.00000e-03*ic_res+1.25000e-01'
+ rm3 = '2.25000e-03*ic_res+4.70000e-02'
+ rm4 = '2.25000e-03*ic_res+4.70000e-02'
+ rm5 = '-2.16840e-19*ic_res*ic_res+1.82500e-03*ic_res+2.85000e-02'
+ rnw = '1.15000e+02*ic_res+1.70000e+03'
+ rp1 = '5.00000e-02*ic_res_poly*ic_res_poly+1.70000e+00*ic_res_poly+4.82000e+01'
+ tol_li = '-5.00000e-09*ic_res'
+ tol_m1 = '-6.25000e-09*ic_res'
+ tol_m2 = '-6.25000e-09*ic_res'
+ tol_m3 = '-1.62500e-08*ic_res'
+ tol_m4 = '-1.62500e-08*ic_res'
+ tol_m5 = '-4.25000e-08*ic_res'
+ tol_nfom = '-1.72500e-08*ic_res'
+ tol_nw = '-1.72500e-08*ic_res'
+ tol_pfom = '-1.50000e-08*ic_res'
+ tol_poly = '-1.02500e-08*ic_res'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield__cor = '3.30000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1__cor = '3.30000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor = '3.62500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3__cor = '2.87500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield__cor = '5.35000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3__cor = '-4.37500e-04*ic_cap*ic_cap+3.25000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield__cor = '5.10000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor = '5.10000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1__cor = '5.62500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor = '4.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor = '4.32500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1__cor = '4.32500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4__cor = '5.20000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1__cor = '4.75000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3__cor = '3.85000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__model__cap_vpp_finger__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield_base__cor = '5.00000e-02*ic_cap+1.00000e+00'

*----------------------------------------------------------
* Include all device model files
*----------------------------------------------------------
* SRAM MOSFETs
*----------------------------------------------------------
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_flash.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_latch.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_pfet_pass.pm3.spice"
*----------------------------------------------------------
* SONOS
*----------------------------------------------------------
.include "../sonos_e/begin_of_life.pm3.spice"
.include "../sonos_p/begin_of_life.pm3.spice"
*----------------------------------------------------------
* Vertical parallel plate (VPP) capacitors
*----------------------------------------------------------
.include "../rescap/sky130_fd_pr__model__cap_vpp_only_mos.model.spice"
.include "../rescap/sky130_fd_pr__model__cap_vpp_only_p.model.spice"
.include "../rescap/sky130_fd_pr__model__cap_vpp_only_pq.model.spice"
*----------------------------------------------------------
* RF MOSFET models
*----------------------------------------------------------
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_mvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"
*----------------------------------------------------------
* Medium-Vt pFET model
*----------------------------------------------------------
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_mvt.pm3.spice"
*----------------------------------------------------------
* Additional resistor models
*----------------------------------------------------------
.include "../rescap/sky130_fd_pr__model__res.model.spice"
