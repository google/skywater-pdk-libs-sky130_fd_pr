* SKY130 legacy discrete models
* Parameters used by res_generic_nd/pd__hv
.param
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = 1.0559e+0
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = 1.0542e+0
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = 1.1193e+0
+ sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult = 1.1801e+0

.include "../../../cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__ss.corner.spice"
