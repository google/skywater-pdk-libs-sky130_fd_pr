* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./parameters_fet_ss.spice created from ./parameters.spice
*
.param sw_tox_lv_corner = {4.148e-09+corner_factor*1.5199999999999948e-10}
.param sw_tox_hv_corner = {1.16e-08+corner_factor*5.000000000000012e-10}
.param sw_polycd = {0.0+corner_factor*5.5e-09} + process_mc_factor*MC_PR_SWITCH*AGAUSS(0,1.5e-09,1)
.param sw_activecd = {0.0+corner_factor*2.25e-08} + process_mc_factor*MC_PR_SWITCH*AGAUSS(0,5e-09,1)
.param sw_nw_rs_mult = {1.0+corner_factor*0.30000000000000004} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.12,1))
.param sw_sky130_fd_pr__pfet_01v8_de_rd_mult = {1.0+corner_factor*0.30000000000000004}
.param sw_nsd_pw_cj = {0.00135+corner_factor*0.00019999999999999987} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_psd_nw_cj = {0.0007408+corner_factor*4.629999999999999e-05} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_nw_pw_cj = {9e-05+corner_factor*1.1999999999999994e-05} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_pw_dnw_cj = {0.0003824+corner_factor*8.069999999999996e-05} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_dnw_sub_cj = {7.743e-05+corner_factor*1.4780000000000004e-05} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_nldd = {1.0+corner_factor*0.19999999999999996} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_vth0_sky130_fd_pr__nfet_01v8 = {0.0+corner_factor*0.015}
.param sw_u0_sky130_fd_pr__nfet_01v8 = {1.0+corner_factor*-0.020000000000000018}
.param sw_vsat_sky130_fd_pr__nfet_01v8 = {1.0+corner_factor*-0.09999999999999998}
.param sw_vth0_sky130_fd_pr__nfet_01v8_lvt = {0.0+corner_factor*0.019}
.param sw_u0_sky130_fd_pr__nfet_01v8_lvt = {1.0+corner_factor*-0.030000000000000027}
.param sw_vth0_sky130_fd_pr__nfet_g5v0d10v5 = {0.0+corner_factor*0.02}
.param sw_u0_sky130_fd_pr__nfet_g5v0d10v5 = {1.0+corner_factor*-0.030000000000000027}
.param sw_vsat_sky130_fd_pr__nfet_g5v0d10v5 = {1.0+corner_factor*-0.09999999999999998}
.param sw_vth0_sky130_fd_pr__nfet_01v8_nat = {0.0+corner_factor*0.02}
.param sw_u0_sky130_fd_pr__nfet_01v8_nat = {1.0+corner_factor*-0.030000000000000027}
.param sw_vth0_sky130_fd_pr__nfet_01v8_zvt = {0.0+corner_factor*0.02} + process_mc_factor*MC_PR_SWITCH*AGAUSS(0,0.007,1)
.param sw_u0_sky130_fd_pr__nfet_01v8_zvt = {1.0+corner_factor*-0.030000000000000027}
.param sw_vth0_sky130_fd_pr__nfet_g5v0d16v0 = {0.0+corner_factor*0.08}
.param sw_u0_sky130_fd_pr__nfet_g5v0d16v0 = {1.0+corner_factor*-0.09999999999999998}
.param sw_vsat_sky130_fd_pr__nfet_g5v0d16v0 = {1.0+corner_factor*-0.25}
.param sw_vth0_sky130_fd_pr__pfet_01v8 = {0.0+corner_factor*-0.01}
.param sw_u0_sky130_fd_pr__pfet_01v8 = {1.0+corner_factor*-0.050000000000000044}
.param sw_vsat_sky130_fd_pr__pfet_01v8 = {1.0+corner_factor*-0.15000000000000002}
.param sw_vth0_sky130_fd_pr__pfet_01v8_lvt = {0.0+corner_factor*-0.09}
.param sw_u0_sky130_fd_pr__pfet_01v8_lvt = {1.0+corner_factor*-0.06999999999999995}
.param sw_vth0_sky130_fd_pr__pfet_01v8_hvt = {0.0+corner_factor*-0.02}
.param sw_u0_sky130_fd_pr__pfet_01v8_hvt = {1.0+corner_factor*-0.06999999999999995}
.param sw_vsat_sky130_fd_pr__pfet_01v8_hvt = {1.0+corner_factor*-0.19999999999999996}
.param sw_vth0_nat_v5 = {-0.0105+corner_factor*0.02441}
.param sw_vth0_sky130_fd_pr__pfet_g5v0d10v5 = {0.0+corner_factor*-0.04}
.param sw_u0_sky130_fd_pr__pfet_g5v0d10v5 = {1.0+corner_factor*-0.06999999999999995}
.param sw_vsat_sky130_fd_pr__pfet_g5v0d10v5 = {1.0+corner_factor*-0.09999999999999998}
.param sw_vth0_sky130_fd_pr__pfet_g5v0d16v0 = {0.0+corner_factor*-0.07}
.param sw_u0_sky130_fd_pr__pfet_g5v0d16v0 = {1.0+corner_factor*-0.06999999999999995}
.param sw_vsat_sky130_fd_pr__pfet_g5v0d16v0 = {1.0+corner_factor*-0.09999999999999998}
