* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
*.PININFO DRAIN:? GATE:? SOURCE:? SUBSTRATE:?
M1 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M2 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M3 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M4 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M5 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M6 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M7 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M8 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M9 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M10 DRAIN GATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M11 SUBSTRATE SUBSTRATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
M12 SUBSTRATE SUBSTRATE SUBSTRATE model_use_only w=7.09 l=0.5 m=1
.ENDS sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50
