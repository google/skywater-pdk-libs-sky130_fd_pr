* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_pfet_01v8_hvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_01v8_hvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_01v8_hvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__special_pfet_01v8_hvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__special_pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__special_pfet_01v8_hvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__special_pfet_01v8_hvt d g s b sky130_fd_pr__special_pfet_01v8_hvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__special_pfet_01v8_hvt__model.0 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.59e-07 wmax = 3.61e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__special_pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = {4.23e-09*sky130_fd_pr__special_pfet_01v8_hvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*sky130_fd_pr__special_pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__special_pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__special_pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__special_pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__special_pfet_01v8_hvt__lint_diff}
*(mismatch parameter sky130_fd_pr__special_pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = {-1.0751186382512+sky130_fd_pr__special_pfet_01v8_hvt__vth0_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__special_pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.915817576187918
+ k2 = {-0.191354581465138+sky130_fd_pr__special_pfet_01v8_hvt__k2_diff_0}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.632029034401906
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__special_pfet_01v8_hvt__voff_slope_spectre)
+ voff = {-0.252068561266462+sky130_fd_pr__special_pfet_01v8_hvt__voff_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__special_pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__special_pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = {3.06838122728761+sky130_fd_pr__special_pfet_01v8_hvt__nfactor_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__special_pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.709002668530266+sky130_fd_pr__special_pfet_01v8_hvt__eta0_diff_0}
+ etab = 0.0119734813782515
+ u0 = {0.00388572612584648+sky130_fd_pr__special_pfet_01v8_hvt__u0_diff_0}
+ ua = {-2.00244775464247e-09+sky130_fd_pr__special_pfet_01v8_hvt__ua_diff_0}
+ ub = {1.8126637343077e-18+sky130_fd_pr__special_pfet_01v8_hvt__ub_diff_0}
+ uc = -3.29420596540557e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {123538.047249085+sky130_fd_pr__special_pfet_01v8_hvt__vsat_diff_0}
+ a0 = {0.999069843161314+sky130_fd_pr__special_pfet_01v8_hvt__a0_diff_0}
+ ags = {1.24999999958161+sky130_fd_pr__special_pfet_01v8_hvt__ags_diff_0}
+ a1 = 0.0
+ a2 = 0.402340703539025
+ b0 = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__b0_diff_0}
+ b1 = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__b1_diff_0}
+ keta = {-0.059104614991198+sky130_fd_pr__special_pfet_01v8_hvt__keta_diff_0}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.626485556768748+sky130_fd_pr__special_pfet_01v8_hvt__pclm_diff_0}
+ pdiblc1 = 0.156960184691247
+ pdiblc2 = 0.00484688249504905
+ pdiblcb = -0.816101282025912
+ drout = 0.999999999574636
+ pscbe1 = 813825374.586324
+ pscbe2 = 9.67821053778591e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__pditsd_diff_0}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__special_pfet_01v8_hvt__rdsw_diff_0}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.66184153982975
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__agidl_diff_0}
+ bgidl = {1000000000.29118+sky130_fd_pr__special_pfet_01v8_hvt__bgidl_diff_0}
+ cgidl = {300.0+sky130_fd_pr__special_pfet_01v8_hvt__cgidl_diff_0}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__special_pfet_01v8_hvt__dlc_diff+sky130_fd_pr__special_pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__special_pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__special_pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__special_pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__special_pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__special_pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__special_pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__special_pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.486150550825388+sky130_fd_pr__special_pfet_01v8_hvt__kt1_diff_0}
+ kt2 = -0.0168844133026869
+ at = 23782.3869663337
+ ute = -0.163199999725863
+ ua1 = 9.15790453404767e-10
+ ub1 = -6.16621741789699e-19
+ uc1 = -1.12531129150376e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__special_pfet_01v8_hvt__tvoff_diff_0}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.ends sky130_fd_pr__special_pfet_01v8_hvt
