* SKY130 Spice File.
.include "../all.spice"
.include "rf.spice"
