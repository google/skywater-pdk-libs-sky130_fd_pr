* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_pr__rf_nfet_20v0_zvt_withptap D PSUB S
X0 D a_n1600_n800# S PSUB sky130_fd_pr__nfet_20v0_nvt w=1.5e+07u l=2.1e+07u
X1 D a_n1600_n800# S PSUB sky130_fd_pr__nfet_20v0_nvt w=1.5e+07u l=2.1e+07u
.ends
