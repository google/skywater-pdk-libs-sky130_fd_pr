* SKY130 Spice File.
*  P+ Poly Preres Corner Parameters
.param
+ sky130_fd_pr__res_high_po__var_mult = -5.0
+ camimc=  1.778e-15  $ Units: farad/micrometer^2
+ cpmimc = 0.03e-15 $ Units: farad/micrometer
+ cvpp_cor = 0.862
+ cvpp3_cor = 0.7
+ cvpp4_cor = 0.7
+ cvpp5_cor = 0.7
+ cm3m2_vpp = 0.446
+ c0m5m4_vpp = 0.804
+ c1m5m4_vpp = 0.766
+ c0m5m4_vpp0p4shield = 0.6046
+ c1m5m4_vpp0p4shield = 0.766
+ c0m4m3_vpp = 0.804
+ c1m4m3_vpp = 0.766
+ c0m5m3_vpp = 0.803
+ c1m5m3_vpp = 0.774
+ cpl2s_vpp = 0.760
+ cpl2s_vpp0p4shield = 0.7511
+ cli2s_vpp = 0.794
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1__cor = 0.810
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1__cor = 0.775
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor = 0.855
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor = 0.827
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield__cor = 0.796
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield__cor = 0.868
+ sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield__cor = 0.786
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1__cor = 0.827
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor = 0.796
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1__cor = 0.868
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3__cor = 0.846
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor = 0.816
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3__cor = 0.885
+ sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3__cor = 0.863
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5__cor = 0.856
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor = 0.856
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor = 0.856
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4__cor = 0.792
+ sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor = 0.8
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4__cor = 0.8
+ sky130_fd_pr__model__cap_vpp_finger__cor = 0.8
+ sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield_base__cor = 0.8
*.param cm3m2_vpp = 0.723
