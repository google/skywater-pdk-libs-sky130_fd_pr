# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__res_high_po_5p73__example1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__res_high_po_5p73__example1 ;
  ORIGIN  2.080000  0.000000 ;
  SIZE  9.890000 BY  5.730000 ;
  OBS
    LAYER li1 ;
      RECT -2.080000 0.000000 0.060000 0.240000 ;
      RECT -2.080000 0.240000 0.080000 5.490000 ;
      RECT -2.080000 5.490000 0.060000 5.730000 ;
      RECT  5.650000 0.240000 7.810000 5.490000 ;
      RECT  5.670000 0.000000 7.810000 0.240000 ;
      RECT  5.670000 5.490000 7.810000 5.730000 ;
    LAYER mcon ;
      RECT -1.970000 0.260000 0.000000 5.470000 ;
      RECT  5.730000 0.260000 7.700000 5.470000 ;
    LAYER met1 ;
      RECT -2.030000 0.200000 0.060000 5.530000 ;
      RECT  5.670000 0.200000 7.760000 5.530000 ;
  END
END sky130_fd_pr__res_high_po_5p73__example1
END LIBRARY
