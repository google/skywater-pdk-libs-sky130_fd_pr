# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_sh_auvia__example_182062124
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_sh_auvia__example_182062124 ;
  ORIGIN  1.790000  2.565000 ;
  SIZE  3.580000 BY  5.130000 ;
  OBS
    LAYER met3 ;
      RECT -1.790000 -2.565000 1.790000 2.565000 ;
    LAYER met4 ;
      RECT -1.790000 -2.565000 1.790000 2.565000 ;
    LAYER via3 ;
      RECT -1.760000 -2.560000 1.760000 2.560000 ;
  END
END sky130_fd_pr__rf_sh_auvia__example_182062124
END LIBRARY
