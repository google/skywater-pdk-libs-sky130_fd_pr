* SKY130 legacy discrete models
* Parameters used by res_generic_nd/pd__hv
.param
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = 9.5405e-1
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = 9.6374e-1
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = 8.7078e-1
+ sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult = 8.4883e-1

.include "../../../cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__ff.corner.spice"
