# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__model__nfet__example1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__model__nfet__example1 ;
  ORIGIN  0.625000  0.130000 ;
  SIZE  1.040000 BY  0.680000 ;
  OBS
    LAYER li1 ;
      RECT -0.565000 -0.020000 -0.055000 0.310000 ;
      RECT  0.205000 -0.020000  0.375000 0.310000 ;
    LAYER mcon ;
      RECT -0.225000 -0.020000 -0.055000 0.150000 ;
    LAYER met1 ;
      RECT -0.255000 -0.080000 -0.025000 0.210000 ;
  END
END sky130_fd_pr__model__nfet__example1
END LIBRARY
