* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param   tc1rsn_h= 1.405e-3
.param   tc2rsn_h= 4.233e-7
.param   tc1rsp_h= 1.369e-3
.param   tc2rsp_h= 1.476e-6

.model sky130_fd_pr__res_generic_nd__hv r tc1r = {tc1rsn_h} tc2r = {tc2rsn_h} rsh = {rdn_hv} dw = {"-tol_nfom/2-nfom_dw/2"} tnom = 30.0
.model sky130_fd_pr__res_generic_pd__hv r tc1r = {tc1rsp_h} tc2r = {tc2rsp_h} rsh = {rdp_hv} dw = {"-tol_pfom/2-pfom_dw/2"} tnom = 30.0

* Resistor model "short" defined with a fixed resistance of 0.01 ohms.
.model short r r=0.01
* If "short" is called as a subcircuit, then this needs to be supported, too.
.subckt short 1 2 SUB l=0 w=0
R0 1 2 short
.ends

* Subcircuit definition HV diffusion resistors

.subckt sky130_fd_pr__res_generic_nd__hv t1 t2 b w=1 l=1
r0 t1 t2 sky130_fd_pr__res_generic_nd__hv w = {w} l = {l}
d0 b t1 sky130_fd_pr__diode_pw2nd_11v0 area='w*l*0.5' pj='w+l'
d1 b t2 sky130_fd_pr__diode_pw2nd_11v0 area='w*l*0.5' pj='w+l'
.ends sky130_fd_pr__res_generic_nd__hv

.subckt sky130_fd_pr__res_generic_pd__hv t1 t2 b w=1 l=1
r0 t1 t2 sky130_fd_pr__res_generic_pd__hv w = {w} l = {l}
d0 t1 b sky130_fd_pr__diode_pd2nw_11v0 area='w*l*0.5' pj='w+l'
d1 t1 b sky130_fd_pr__diode_pd2nw_11v0 area='w*l*0.5' pj='w+l'
.ends sky130_fd_pr__res_generic_pd__hv

* Simple subcircuit definitions for legacy fixed-width resistors

.subckt sky130_fd_pr__res_high_po_0p35 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_high_po l=l w=0.35 mult=mult
.ends sky130_fd_pr__res_high_po_0p35

.subckt sky130_fd_pr__res_high_po_0p69 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_high_po l=l w=0.69 mult=mult
.ends sky130_fd_pr__res_high_po_0p69

.subckt sky130_fd_pr__res_high_po_1p41 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_high_po l=l w=1.41 mult=mult
.ends sky130_fd_pr__res_high_po_1p41

.subckt sky130_fd_pr__res_high_po_2p85 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_high_po l=l w=2.85 mult=mult
.ends sky130_fd_pr__res_high_po_2p85

.subckt sky130_fd_pr__res_high_po_5p73 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_high_po l=l w=5.73 mult=mult
.ends sky130_fd_pr__res_high_po_5p73

.subckt sky130_fd_pr__res_xhigh_po_0p35 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_xhigh_po l=l w=0.35 mult=mult
.ends sky130_fd_pr__res_xhigh_po_0p35

.subckt sky130_fd_pr__res_xhigh_po_0p69 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_xhigh_po l=l w=0.69 mult=mult
.ends sky130_fd_pr__res_xhigh_po_0p69

.subckt sky130_fd_pr__res_xhigh_po_1p41 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_xhigh_po l=l w=1.41 mult=mult
.ends sky130_fd_pr__res_xhigh_po_1p41

.subckt sky130_fd_pr__res_xhigh_po_2p85 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_xhigh_po l=l w=2.85 mult=mult
.ends sky130_fd_pr__res_xhigh_po_2p85

.subckt sky130_fd_pr__res_xhigh_po_5p73 r0 r1 sub mult=1 l=1
x0 r0 r1 sub sky130_fd_pr__res_xhigh_po l=l w=5.73 mult=mult
.ends sky130_fd_pr__res_xhigh_po_5p73
