# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__via_m2m3__example4
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__via_m2m3__example4 ;
  ORIGIN  0.025000  0.000000 ;
  SIZE  0.330000 BY  0.370000 ;
  OBS
    LAYER met2 ;
      RECT 0.000000 0.000000 0.280000 0.370000 ;
    LAYER met3 ;
      RECT -0.025000 0.020000 0.305000 0.350000 ;
    LAYER via2 ;
      RECT 0.000000 0.045000 0.280000 0.325000 ;
  END
END sky130_fd_pr__via_m2m3__example4
END LIBRARY
