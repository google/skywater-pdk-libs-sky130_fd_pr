# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__genrivetdlring__example_179576876
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__genrivetdlring__example_179576876 ;
  ORIGIN  0.190000  0.190000 ;
  SIZE  65.16000 BY  65.16000 ;
  OBS
    LAYER met4 ;
      RECT -0.190000  6.235000  0.990000  7.415000 ;
      RECT -0.190000  7.835000  0.990000  9.015000 ;
      RECT -0.190000  9.435000  0.990000 10.615000 ;
      RECT -0.190000 11.035000  0.990000 12.215000 ;
      RECT -0.190000 12.635000  0.990000 13.815000 ;
      RECT -0.190000 14.235000  0.990000 15.415000 ;
      RECT -0.190000 15.835000  0.990000 17.015000 ;
      RECT -0.190000 17.435000  0.990000 18.615000 ;
      RECT -0.190000 19.035000  0.990000 20.215000 ;
      RECT -0.190000 20.635000  0.990000 21.815000 ;
      RECT -0.190000 22.235000  0.990000 23.415000 ;
      RECT -0.190000 23.835000  0.990000 25.015000 ;
      RECT -0.190000 25.435000  0.990000 26.615000 ;
      RECT -0.190000 27.035000  0.990000 28.215000 ;
      RECT -0.190000 28.635000  0.990000 29.815000 ;
      RECT -0.190000 30.235000  0.990000 31.415000 ;
      RECT -0.190000 31.835000  0.990000 33.015000 ;
      RECT -0.190000 33.435000  0.990000 34.615000 ;
      RECT -0.190000 35.035000  0.990000 36.215000 ;
      RECT -0.190000 36.635000  0.990000 37.815000 ;
      RECT -0.190000 38.235000  0.990000 39.415000 ;
      RECT -0.190000 39.835000  0.990000 41.015000 ;
      RECT -0.190000 41.435000  0.990000 42.615000 ;
      RECT -0.190000 43.035000  0.990000 44.215000 ;
      RECT -0.190000 44.635000  0.990000 45.815000 ;
      RECT -0.190000 46.235000  0.990000 47.415000 ;
      RECT -0.190000 47.835000  0.990000 49.015000 ;
      RECT -0.190000 49.435000  0.990000 50.615000 ;
      RECT -0.190000 51.035000  0.990000 52.215000 ;
      RECT -0.190000 52.635000  0.990000 53.815000 ;
      RECT -0.190000 54.235000  0.990000 55.415000 ;
      RECT -0.190000 55.835000  0.990000 57.015000 ;
      RECT -0.190000 57.435000  0.990000 58.615000 ;
      RECT  1.355000  4.620000  2.535000  5.800000 ;
      RECT  1.425000 59.050000  2.605000 60.230000 ;
      RECT  2.955000  3.020000  4.135000  4.200000 ;
      RECT  3.025000 60.650000  4.205000 61.830000 ;
      RECT  4.555000  1.420000  5.735000  2.600000 ;
      RECT  4.625000 62.250000  5.805000 63.430000 ;
      RECT  6.165000 -0.190000  7.345000  0.990000 ;
      RECT  6.235000 63.790000  7.415000 64.970000 ;
      RECT  7.765000 -0.190000  8.945000  0.990000 ;
      RECT  7.835000 63.790000  9.015000 64.970000 ;
      RECT  9.365000 -0.190000 10.545000  0.990000 ;
      RECT  9.435000 63.790000 10.615000 64.970000 ;
      RECT 10.965000 -0.190000 12.145000  0.990000 ;
      RECT 11.035000 63.790000 12.215000 64.970000 ;
      RECT 12.565000 -0.190000 13.745000  0.990000 ;
      RECT 12.635000 63.790000 13.815000 64.970000 ;
      RECT 14.165000 -0.190000 15.345000  0.990000 ;
      RECT 14.235000 63.790000 15.415000 64.970000 ;
      RECT 15.765000 -0.190000 16.945000  0.990000 ;
      RECT 15.835000 63.790000 17.015000 64.970000 ;
      RECT 17.365000 -0.190000 18.545000  0.990000 ;
      RECT 17.435000 63.790000 18.615000 64.970000 ;
      RECT 18.965000 -0.190000 20.145000  0.990000 ;
      RECT 19.035000 63.790000 20.215000 64.970000 ;
      RECT 20.565000 -0.190000 21.745000  0.990000 ;
      RECT 20.635000 63.790000 21.815000 64.970000 ;
      RECT 22.165000 -0.190000 23.345000  0.990000 ;
      RECT 22.235000 63.790000 23.415000 64.970000 ;
      RECT 23.765000 -0.190000 24.945000  0.990000 ;
      RECT 23.835000 63.790000 25.015000 64.970000 ;
      RECT 25.365000 -0.190000 26.545000  0.990000 ;
      RECT 25.435000 63.790000 26.615000 64.970000 ;
      RECT 26.965000 -0.190000 28.145000  0.990000 ;
      RECT 27.035000 63.790000 28.215000 64.970000 ;
      RECT 28.565000 -0.190000 29.745000  0.990000 ;
      RECT 28.635000 63.790000 29.815000 64.970000 ;
      RECT 30.165000 -0.190000 31.345000  0.990000 ;
      RECT 30.235000 63.790000 31.415000 64.970000 ;
      RECT 31.765000 -0.190000 32.945000  0.990000 ;
      RECT 31.835000 63.790000 33.015000 64.970000 ;
      RECT 33.365000 -0.190000 34.545000  0.990000 ;
      RECT 33.435000 63.790000 34.615000 64.970000 ;
      RECT 34.965000 -0.190000 36.145000  0.990000 ;
      RECT 35.035000 63.790000 36.215000 64.970000 ;
      RECT 36.565000 -0.190000 37.745000  0.990000 ;
      RECT 36.635000 63.790000 37.815000 64.970000 ;
      RECT 38.165000 -0.190000 39.345000  0.990000 ;
      RECT 38.235000 63.790000 39.415000 64.970000 ;
      RECT 39.765000 -0.190000 40.945000  0.990000 ;
      RECT 39.835000 63.790000 41.015000 64.970000 ;
      RECT 41.365000 -0.190000 42.545000  0.990000 ;
      RECT 41.435000 63.790000 42.615000 64.970000 ;
      RECT 42.965000 -0.190000 44.145000  0.990000 ;
      RECT 43.035000 63.790000 44.215000 64.970000 ;
      RECT 44.565000 -0.190000 45.745000  0.990000 ;
      RECT 44.635000 63.790000 45.815000 64.970000 ;
      RECT 46.165000 -0.190000 47.345000  0.990000 ;
      RECT 46.235000 63.790000 47.415000 64.970000 ;
      RECT 47.765000 -0.190000 48.945000  0.990000 ;
      RECT 47.835000 63.790000 49.015000 64.970000 ;
      RECT 49.365000 -0.190000 50.545000  0.990000 ;
      RECT 49.435000 63.790000 50.615000 64.970000 ;
      RECT 50.965000 -0.190000 52.145000  0.990000 ;
      RECT 51.035000 63.790000 52.215000 64.970000 ;
      RECT 52.565000 -0.190000 53.745000  0.990000 ;
      RECT 52.635000 63.790000 53.815000 64.970000 ;
      RECT 54.165000 -0.190000 55.345000  0.990000 ;
      RECT 54.235000 63.790000 55.415000 64.970000 ;
      RECT 55.765000 -0.190000 56.945000  0.990000 ;
      RECT 55.835000 63.790000 57.015000 64.970000 ;
      RECT 57.365000 -0.190000 58.545000  0.990000 ;
      RECT 57.435000 63.790000 58.615000 64.970000 ;
      RECT 58.975000  1.350000 60.155000  2.530000 ;
      RECT 59.045000 62.180000 60.225000 63.360000 ;
      RECT 60.575000  2.950000 61.755000  4.130000 ;
      RECT 60.645000 60.580000 61.825000 61.760000 ;
      RECT 62.175000  4.550000 63.355000  5.730000 ;
      RECT 62.245000 58.980000 63.425000 60.160000 ;
      RECT 63.790000  6.165000 64.970000  7.345000 ;
      RECT 63.790000  7.765000 64.970000  8.945000 ;
      RECT 63.790000  9.365000 64.970000 10.545000 ;
      RECT 63.790000 10.965000 64.970000 12.145000 ;
      RECT 63.790000 12.565000 64.970000 13.745000 ;
      RECT 63.790000 14.165000 64.970000 15.345000 ;
      RECT 63.790000 15.765000 64.970000 16.945000 ;
      RECT 63.790000 17.365000 64.970000 18.545000 ;
      RECT 63.790000 18.965000 64.970000 20.145000 ;
      RECT 63.790000 20.565000 64.970000 21.745000 ;
      RECT 63.790000 22.165000 64.970000 23.345000 ;
      RECT 63.790000 23.765000 64.970000 24.945000 ;
      RECT 63.790000 25.365000 64.970000 26.545000 ;
      RECT 63.790000 26.965000 64.970000 28.145000 ;
      RECT 63.790000 28.565000 64.970000 29.745000 ;
      RECT 63.790000 30.165000 64.970000 31.345000 ;
      RECT 63.790000 31.765000 64.970000 32.945000 ;
      RECT 63.790000 33.365000 64.970000 34.545000 ;
      RECT 63.790000 34.965000 64.970000 36.145000 ;
      RECT 63.790000 36.565000 64.970000 37.745000 ;
      RECT 63.790000 38.165000 64.970000 39.345000 ;
      RECT 63.790000 39.765000 64.970000 40.945000 ;
      RECT 63.790000 41.365000 64.970000 42.545000 ;
      RECT 63.790000 42.965000 64.970000 44.145000 ;
      RECT 63.790000 44.565000 64.970000 45.745000 ;
      RECT 63.790000 46.165000 64.970000 47.345000 ;
      RECT 63.790000 47.765000 64.970000 48.945000 ;
      RECT 63.790000 49.365000 64.970000 50.545000 ;
      RECT 63.790000 50.965000 64.970000 52.145000 ;
      RECT 63.790000 52.565000 64.970000 53.745000 ;
      RECT 63.790000 54.165000 64.970000 55.345000 ;
      RECT 63.790000 55.765000 64.970000 56.945000 ;
      RECT 63.790000 57.365000 64.970000 58.545000 ;
    LAYER met5 ;
      RECT -0.190000  6.235000  0.990000  7.415000 ;
      RECT -0.190000  7.835000  0.990000  9.015000 ;
      RECT -0.190000  9.435000  0.990000 10.615000 ;
      RECT -0.190000 11.035000  0.990000 12.215000 ;
      RECT -0.190000 12.635000  0.990000 13.815000 ;
      RECT -0.190000 14.235000  0.990000 15.415000 ;
      RECT -0.190000 15.835000  0.990000 17.015000 ;
      RECT -0.190000 17.435000  0.990000 18.615000 ;
      RECT -0.190000 19.035000  0.990000 20.215000 ;
      RECT -0.190000 20.635000  0.990000 21.815000 ;
      RECT -0.190000 22.235000  0.990000 23.415000 ;
      RECT -0.190000 23.835000  0.990000 25.015000 ;
      RECT -0.190000 25.435000  0.990000 26.615000 ;
      RECT -0.190000 27.035000  0.990000 28.215000 ;
      RECT -0.190000 28.635000  0.990000 29.815000 ;
      RECT -0.190000 30.235000  0.990000 31.415000 ;
      RECT -0.190000 31.835000  0.990000 33.015000 ;
      RECT -0.190000 33.435000  0.990000 34.615000 ;
      RECT -0.190000 35.035000  0.990000 36.215000 ;
      RECT -0.190000 36.635000  0.990000 37.815000 ;
      RECT -0.190000 38.235000  0.990000 39.415000 ;
      RECT -0.190000 39.835000  0.990000 41.015000 ;
      RECT -0.190000 41.435000  0.990000 42.615000 ;
      RECT -0.190000 43.035000  0.990000 44.215000 ;
      RECT -0.190000 44.635000  0.990000 45.815000 ;
      RECT -0.190000 46.235000  0.990000 47.415000 ;
      RECT -0.190000 47.835000  0.990000 49.015000 ;
      RECT -0.190000 49.435000  0.990000 50.615000 ;
      RECT -0.190000 51.035000  0.990000 52.215000 ;
      RECT -0.190000 52.635000  0.990000 53.815000 ;
      RECT -0.190000 54.235000  0.990000 55.415000 ;
      RECT -0.190000 55.835000  0.990000 57.015000 ;
      RECT -0.190000 57.435000  0.990000 58.615000 ;
      RECT  1.355000  4.620000  2.535000  5.800000 ;
      RECT  1.425000 59.050000  2.605000 60.230000 ;
      RECT  2.955000  3.020000  4.135000  4.200000 ;
      RECT  3.025000 60.650000  4.205000 61.830000 ;
      RECT  4.555000  1.420000  5.735000  2.600000 ;
      RECT  4.625000 62.250000  5.805000 63.430000 ;
      RECT  6.165000 -0.190000  7.345000  0.990000 ;
      RECT  6.235000 63.790000  7.415000 64.970000 ;
      RECT  7.765000 -0.190000  8.945000  0.990000 ;
      RECT  7.835000 63.790000  9.015000 64.970000 ;
      RECT  9.365000 -0.190000 10.545000  0.990000 ;
      RECT  9.435000 63.790000 10.615000 64.970000 ;
      RECT 10.965000 -0.190000 12.145000  0.990000 ;
      RECT 11.035000 63.790000 12.215000 64.970000 ;
      RECT 12.565000 -0.190000 13.745000  0.990000 ;
      RECT 12.635000 63.790000 13.815000 64.970000 ;
      RECT 14.165000 -0.190000 15.345000  0.990000 ;
      RECT 14.235000 63.790000 15.415000 64.970000 ;
      RECT 15.765000 -0.190000 16.945000  0.990000 ;
      RECT 15.835000 63.790000 17.015000 64.970000 ;
      RECT 17.365000 -0.190000 18.545000  0.990000 ;
      RECT 17.435000 63.790000 18.615000 64.970000 ;
      RECT 18.965000 -0.190000 20.145000  0.990000 ;
      RECT 19.035000 63.790000 20.215000 64.970000 ;
      RECT 20.565000 -0.190000 21.745000  0.990000 ;
      RECT 20.635000 63.790000 21.815000 64.970000 ;
      RECT 22.165000 -0.190000 23.345000  0.990000 ;
      RECT 22.235000 63.790000 23.415000 64.970000 ;
      RECT 23.765000 -0.190000 24.945000  0.990000 ;
      RECT 23.835000 63.790000 25.015000 64.970000 ;
      RECT 25.365000 -0.190000 26.545000  0.990000 ;
      RECT 25.435000 63.790000 26.615000 64.970000 ;
      RECT 26.965000 -0.190000 28.145000  0.990000 ;
      RECT 27.035000 63.790000 28.215000 64.970000 ;
      RECT 28.565000 -0.190000 29.745000  0.990000 ;
      RECT 28.635000 63.790000 29.815000 64.970000 ;
      RECT 30.165000 -0.190000 31.345000  0.990000 ;
      RECT 30.235000 63.790000 31.415000 64.970000 ;
      RECT 31.765000 -0.190000 32.945000  0.990000 ;
      RECT 31.835000 63.790000 33.015000 64.970000 ;
      RECT 33.365000 -0.190000 34.545000  0.990000 ;
      RECT 33.435000 63.790000 34.615000 64.970000 ;
      RECT 34.965000 -0.190000 36.145000  0.990000 ;
      RECT 35.035000 63.790000 36.215000 64.970000 ;
      RECT 36.565000 -0.190000 37.745000  0.990000 ;
      RECT 36.635000 63.790000 37.815000 64.970000 ;
      RECT 38.165000 -0.190000 39.345000  0.990000 ;
      RECT 38.235000 63.790000 39.415000 64.970000 ;
      RECT 39.765000 -0.190000 40.945000  0.990000 ;
      RECT 39.835000 63.790000 41.015000 64.970000 ;
      RECT 41.365000 -0.190000 42.545000  0.990000 ;
      RECT 41.435000 63.790000 42.615000 64.970000 ;
      RECT 42.965000 -0.190000 44.145000  0.990000 ;
      RECT 43.035000 63.790000 44.215000 64.970000 ;
      RECT 44.565000 -0.190000 45.745000  0.990000 ;
      RECT 44.635000 63.790000 45.815000 64.970000 ;
      RECT 46.165000 -0.190000 47.345000  0.990000 ;
      RECT 46.235000 63.790000 47.415000 64.970000 ;
      RECT 47.765000 -0.190000 48.945000  0.990000 ;
      RECT 47.835000 63.790000 49.015000 64.970000 ;
      RECT 49.365000 -0.190000 50.545000  0.990000 ;
      RECT 49.435000 63.790000 50.615000 64.970000 ;
      RECT 50.965000 -0.190000 52.145000  0.990000 ;
      RECT 51.035000 63.790000 52.215000 64.970000 ;
      RECT 52.565000 -0.190000 53.745000  0.990000 ;
      RECT 52.635000 63.790000 53.815000 64.970000 ;
      RECT 54.165000 -0.190000 55.345000  0.990000 ;
      RECT 54.235000 63.790000 55.415000 64.970000 ;
      RECT 55.765000 -0.190000 56.945000  0.990000 ;
      RECT 55.835000 63.790000 57.015000 64.970000 ;
      RECT 57.365000 -0.190000 58.545000  0.990000 ;
      RECT 57.435000 63.790000 58.615000 64.970000 ;
      RECT 58.975000  1.350000 60.155000  2.530000 ;
      RECT 59.045000 62.180000 60.225000 63.360000 ;
      RECT 60.575000  2.950000 61.755000  4.130000 ;
      RECT 60.645000 60.580000 61.825000 61.760000 ;
      RECT 62.175000  4.550000 63.355000  5.730000 ;
      RECT 62.245000 58.980000 63.425000 60.160000 ;
      RECT 63.790000  6.165000 64.970000  7.345000 ;
      RECT 63.790000  7.765000 64.970000  8.945000 ;
      RECT 63.790000  9.365000 64.970000 10.545000 ;
      RECT 63.790000 10.965000 64.970000 12.145000 ;
      RECT 63.790000 12.565000 64.970000 13.745000 ;
      RECT 63.790000 14.165000 64.970000 15.345000 ;
      RECT 63.790000 15.765000 64.970000 16.945000 ;
      RECT 63.790000 17.365000 64.970000 18.545000 ;
      RECT 63.790000 18.965000 64.970000 20.145000 ;
      RECT 63.790000 20.565000 64.970000 21.745000 ;
      RECT 63.790000 22.165000 64.970000 23.345000 ;
      RECT 63.790000 23.765000 64.970000 24.945000 ;
      RECT 63.790000 25.365000 64.970000 26.545000 ;
      RECT 63.790000 26.965000 64.970000 28.145000 ;
      RECT 63.790000 28.565000 64.970000 29.745000 ;
      RECT 63.790000 30.165000 64.970000 31.345000 ;
      RECT 63.790000 31.765000 64.970000 32.945000 ;
      RECT 63.790000 33.365000 64.970000 34.545000 ;
      RECT 63.790000 34.965000 64.970000 36.145000 ;
      RECT 63.790000 36.565000 64.970000 37.745000 ;
      RECT 63.790000 38.165000 64.970000 39.345000 ;
      RECT 63.790000 39.765000 64.970000 40.945000 ;
      RECT 63.790000 41.365000 64.970000 42.545000 ;
      RECT 63.790000 42.965000 64.970000 44.145000 ;
      RECT 63.790000 44.565000 64.970000 45.745000 ;
      RECT 63.790000 46.165000 64.970000 47.345000 ;
      RECT 63.790000 47.765000 64.970000 48.945000 ;
      RECT 63.790000 49.365000 64.970000 50.545000 ;
      RECT 63.790000 50.965000 64.970000 52.145000 ;
      RECT 63.790000 52.565000 64.970000 53.745000 ;
      RECT 63.790000 54.165000 64.970000 55.345000 ;
      RECT 63.790000 55.765000 64.970000 56.945000 ;
      RECT 63.790000 57.365000 64.970000 58.545000 ;
  END
END sky130_fd_pr__genrivetdlring__example_179576876
END LIBRARY
