* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
*   mismatch {
*     }
* }
.subckt  sky130_fd_pr__res_high_po_0p35 r0 r1 b
+ 
.param  w = 0.350 l = 5 mult = 1.0
+ 
+ body_pelgrom = 0.0347
+ rend_mm = 0.085
+ rcon = 589.99
+ rsheet = 1112.41
+ tc1_voltco = -7.1e-3
+ vc1_body = -8.46e-3
+ vc2_body = 1.97e-3
+ vc3_body = 3.30e-5
+ vc1_raw_end = -2.02e-2
+ vc2_raw_end = 1.55e-1
+ vc3_raw_end = 4.61e-2
+ r0_var = 50.97
+ r1_var = 34.74
+ vc1_end = {vc1_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))}
+ vc2_end = {vc2_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))}
+ vc3_end = {vc3_raw_end/pwr(l,0.5)*(1+tc1_voltco*(temper-30))}
+ rtot_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2*pow(r0_var,2)+pow((r1_var*l),2))}
+ rend_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2)*r0_var}
+ rbody_var = {rtot_var-rend_var}
+ res_match = {(body_pelgrom/sqrt(w*l*mult))*sky130_fd_pr__res_high_po__slope_spectre}
+ rend = {(rcon+rend_var)*(1+rend_mm/sqrt(mult)*sky130_fd_pr__res_high_po__con_slope_spectre)}
+ rbody = {(l*rsheet+rbody_var)*(1+res_match)}
rend r0 ra r = {rend*(1+min((abs(v(r0,r1))-1.7),0.3)*vc1_end+pow(min(abs(v(r0,r1))-1.7,0.3),2)*vc2_end+pow(min(abs(v(r0,r1))-1.7,0.3),3)*vc3_end)}
rhrpoly_0p35 ra r1 r = {rbody*(1+abs(v(r0,r1))*vc1_body+pow(abs(v(r0,r1)),2)*vc2_body+pow(abs(v(r0,r1)),3)*vc3_body)}
+ tc1 = 0.514e-3
+ tc2 = 0.122e-5
*+ tnom=30
c1 r0 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2}
c2 r1 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2}
.ends sky130_fd_pr__res_high_po_0p35
