* Test the parsers
*---------------------------------------------------------------------
* It should be possible to run both ngspice and Xyce on this simple
* test circuit and have them run without flagging an error.
* This is clearly not exhaustive;  just a quick check on basic syntax
*---------------------------------------------------------------------
.lib sky130.lib.spice tt
Xtest 1 2 3 0 sky130_fd_pr__nfet_01v8 l=2 w=3
.op
.end
