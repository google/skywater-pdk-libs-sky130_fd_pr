* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre = 0.0
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre = 0.0
.param sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre = 0.0
.param sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM02 d g s b sky130_fd_pr__rf_pfet_01v8_bM02__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.0 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.62e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.022+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.784e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0}
+ ua = {-2.45e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_0}
+ ub = {2.075e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_0}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_0}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00307+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_0}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_0}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_0}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2969+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_0+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.23+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_0+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4678
+ pdiblc1 = 0.235
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4527
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.05627
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.556+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_0}
+ kt2 = -0.122
+ at = 4.554e+4
+ ute = -0.39
+ ua1 = 1.346e-10
+ ub1 = 4.516e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {6e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.6e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {2.12e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {-7e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0024*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.0862
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.0
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.1 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.62e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.984+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.217e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1}
+ ua = {-2.37e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_1}
+ ub = {1.99e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_1}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_1}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00305+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_1}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_1}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_1}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3374+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_1+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.99+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_1+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4678
+ pdiblc1 = 7.656e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5264
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0521
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.556+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_1}
+ kt2 = -0.122
+ at = 4.554e+4
+ ute = -0.39
+ ua1 = 1.346e-10
+ ub1 = 4.516e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {7e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.7e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {2.12e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {-2e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0023*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.0862
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.0
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.2 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.62e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.945+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.4e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2}
+ ua = {-2.199e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_2}
+ ub = {1.855e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_2}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_2}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.003331+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_2}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_2}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_2}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3104+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_2+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.87+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_2+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.3036
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4678
+ pdiblc1 = 0.1
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.7475
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0521
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.556+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_2}
+ kt2 = -0.122
+ at = 4.554e+4
+ ute = -0.39
+ ua1 = 1.346e-10
+ ub1 = 4.516e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.4e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {2.12e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {-4e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0023*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.0862
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.0
.ends sky130_fd_pr__rf_pfet_01v8_bM02
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00 d g s b
+ 
.param  l = 1 w = 3.01 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM02W3p00 d g s b sky130_fd_pr__rf_pfet_01v8_bM02__model l = {l} w = 3.01 nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.3 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.2e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3}
+ ua = {-2.307e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_3}
+ ub = {1.975e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_3}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_3}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00431+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_3}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_3}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_3}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3297+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_3+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_3+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.006804
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.279
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.3382
+ pdiblc1 = 0.24
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4851
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.1
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5203+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_3}
+ kt2 = -0.122
+ at = 1.916e+4
+ ute = -0.189
+ ua1 = 1.346e-10
+ ub1 = 9.851e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {8e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.555e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {4.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.52e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {6e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.0
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0024*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.8
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.005+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.2e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4}
+ ua = {-2.197e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_4}
+ ub = {1.859e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_4}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_4}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00429+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_4}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_4}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_4}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_4+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_4+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.006804
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.279
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2949
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4851
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.1
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.52026+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_4}
+ kt2 = -0.122
+ at = 1.916e+4
+ ute = -0.189
+ ua1 = 1.346e-10
+ ub1 = 9.851e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.05e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.455e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {7e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.002*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.8
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.5e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.5 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.976+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.976e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5}
+ ua = {-2.187e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_5}
+ ub = {1.834e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_5}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_5}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00365+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_5}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_5}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_5}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_5+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_5+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0063
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.31
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5899
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5053
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.03747
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.52026+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_5}
+ kt2 = -0.122
+ at = 1.916e+4
+ ute = -0.189
+ ua1 = 1.346e-10
+ ub1 = 9.851e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.2e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.455e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {7e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.ends sky130_fd_pr__rf_pfet_01v8_bM02W3p00
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00 d g s b
+ 
.param  l = 1 w = 5.05 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM02W5p00 d g s b sky130_fd_pr__rf_pfet_01v8_bM02__model l = {l} w = 5.05 nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.6 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.058+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.7e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6}
+ ua = {-2.311e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_6}
+ ub = {1.91e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_6}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_6}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.004327+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_6}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_6}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_6}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_6+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope/sqrt(l*w*mult))}
+ nfactor = {5.651+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_6+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0066
+ cdscb = 0.0
+ cdscd = 0.0039
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.298
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5309
+ pdiblc1 = 0.248
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4188
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.07242
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.56212+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_6}
+ kt2 = -0.122
+ at = 2.705e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {200*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {7.4e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1.3e-08+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.021+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.84e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7}
+ ua = {-2.321e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_7}
+ ub = {1.953e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_7}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_7}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0037+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_7}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_7}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_7}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3074+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_7+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_7+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0046
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4186
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.627
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.05346
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.56212+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_7}
+ kt2 = -0.122
+ at = 3.472e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {200*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.3e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1.4e-08+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM02__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.977+sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.708e+04+sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8}
+ ua = {-2.21e-09+sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_8}
+ ub = {1.824e-18+sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_8}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_8}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00375+sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_8}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_8}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_8}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_8+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_8+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.298
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5899
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5264
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0457
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5162+sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_8}
+ kt2 = -0.122
+ at = 4.321e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {200*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {9.9e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.505e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.ends sky130_fd_pr__rf_pfet_01v8_bM02W5p00
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM04 d g s b sky130_fd_pr__rf_pfet_01v8_bM04__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.0 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.044+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.908e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0}
+ ua = {-2.368e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_0}
+ ub = {1.997e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_0}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_0}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00329+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_0}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_0}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_0}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.345+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_0+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.36+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_0+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.00043
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5085
+ pdiblc1 = 0.12
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.379
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.05667
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_0}
+ kt2 = -0.122
+ at = 3.02e+4
+ ute = -0.036
+ ua1 = 1.992e-10
+ ub1 = 4.398e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {1600*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {8.2e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.7e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.455e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {2.12e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {6e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0015*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.1 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.005+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.808e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1}
+ ua = {-2.325e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_1}
+ ub = {1.939e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_1}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_1}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.003126+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_1}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_1}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_1}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3248+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_1+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_1+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5085
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5264
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0457
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.570+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_1}
+ kt2 = -0.122
+ at = 2.796e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 4.398e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {1600*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {9.2e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.7e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.455e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {2.12e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {6e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0015*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3.2e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.2 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.62e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.955+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.364e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2}
+ ua = {-2.199e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_2}
+ ub = {1.855e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_2}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_2}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.003331+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_2}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_2}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_2}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3104+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_2+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.87+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_2+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1799
+ etab = -0.07835
+ dsub = 0.3036
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4678
+ pdiblc1 = 0.1
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.7475
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0521
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.556+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_2}
+ kt2 = -0.122
+ at = 3.598e+4
+ ute = -0.39
+ ua1 = 1.346e-10
+ ub1 = 4.516e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {1600*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.25e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 2.0e-12
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.3e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.7e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {-4e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.002*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.0862
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.8e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.0
.ends sky130_fd_pr__rf_pfet_01v8_bM04
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00 d g s b
+ 
.param  l = 1 w = 3.01 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM04W3p00 d g s b sky130_fd_pr__rf_pfet_01v8_bM04__model l = {l} w = 3.01 nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.3 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.1e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3}
+ ua = {-2.307e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_3}
+ ub = {1.975e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_3}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_3}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00431+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_3}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_3}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_3}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3297+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_3+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_3+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.006804
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1612
+ etab = -0.07835
+ dsub = 0.279
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.3382
+ pdiblc1 = 0.2448
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4366
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.1
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5515+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_3}
+ kt2 = -0.122
+ at = 2.299e+4
+ ute = -0.1436
+ ua1 = 3.138e-10
+ ub1 = 4.531e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.2e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.1e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.055e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {4.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {6e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.0
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0024*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.8
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.4e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.021+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.912e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4}
+ ua = {-2.219e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_4}
+ ub = {1.915e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_4}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_4}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.004419+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_4}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_4}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_4}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_4+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.242+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_4+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.006804
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.279
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2949
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4851
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.1
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5203+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_4}
+ kt2 = -0.122
+ at = 1.916e+4
+ ute = -0.189
+ ua1 = 1.346e-10
+ ub1 = 9.851e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.25e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.7e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.3e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {7e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.8
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.5 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.983+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.743e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5}
+ ua = {-2.187e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_5}
+ ub = {1.852e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_5}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_5}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00365+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_5}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_5}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_5}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_5+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.531+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_5+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0063
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.31
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5899
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5053
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.03747
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5203+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_5}
+ kt2 = -0.122
+ at = 1.916e+4
+ ute = -0.189
+ ua1 = 1.346e-10
+ ub1 = 9.851e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {800*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.05e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.155e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {7e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.002*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.6e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.ends sky130_fd_pr__rf_pfet_01v8_bM04W3p00
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00 d g s b
+ 
.param  l = 1 w = 5.05 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__rf_pfet_01v8_bM04W5p00 d g s b sky130_fd_pr__rf_pfet_01v8_bM04__model l = {l} w = 5.05 nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.6 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.079+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.7e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6}
+ ua = {-2.311e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_6}
+ ub = {1.948e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_6}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_6}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.004327+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_6}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_6}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_6}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_6+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.103+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_6+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0066
+ cdscb = 0.0
+ cdscd = 0.0039
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.298
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5309
+ pdiblc1 = 0.248
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.4188
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.07242
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5621+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_6}
+ kt2 = -0.122
+ at = 2.705e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {7.4e-07+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.52e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1.3e-08+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0022*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {3e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.026+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {7.213e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7}
+ ua = {-2.328e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_7}
+ ub = {1.953e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_7}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_7}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0037+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_7}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_7}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_7}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3074+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_7+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {6.012+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_7+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0046
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.2663
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.4186
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.627
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.05346
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5621+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_7}
+ kt2 = -0.122
+ at = 3.472e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {0.85e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.5e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1.105e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.72e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1.4e-08+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0017*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.7e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.model sky130_fd_pr__rf_pfet_01v8_bM04__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.399e-08+sky130_fd_pr__rf_pfet_01v8_b__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.304e-09+sky130_fd_pr__rf_pfet_01v8_b__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.786e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 3.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 1.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 2.5e+7
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult+sky130_fd_pr__rf_pfet_01v8__b_toxe_slope_spectre*(4.23e-09*sky130_fd_pr__rf_pfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_pfet_01v8__b_toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.6e+17
+ nsd = 1.0e+20
+ rshg = {49.2+sky130_fd_pr__rf_pfet_01v8_b__rshg_diff}
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9895+sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8+sky130_fd_pr__rf_pfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.038
+ k2 = {-0.1734+sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8}
+ k3 = -15.85
+ dvt0 = 4.585
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.977
+ dvt1w = 1.147e+6
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {6.488e+04+sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8}
+ ua = {-2.21e-09+sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_8}
+ ub = {1.851e-18+sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_8}
+ uc = 2.523e-13
+ rdsw = {547.9+sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_8}
+ prwb = -0.3235
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00375+sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8}
+ a0 = {0.8909+sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_8}
+ keta = 0.0239
+ a1 = 0.0
+ a2 = 0.6419
+ ags = {1.25+sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_8}
+ b0 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_8}
+ b1 = {0+sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 547.9
+ rdwmin = 0.0
+ rsw = 547.9
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.3364+sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_8+sky130_fd_pr__rf_pfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_voff_slope1/sqrt(l*w*mult))}
+ nfactor = {5.892+sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_8+sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope_spectre*(sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1/sqrt(l*w*mult))}
+ cit = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = 0.1874
+ etab = -0.07835
+ dsub = 0.298
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.5899
+ pdiblc1 = 4.4e-11
+ pdiblc2 = 0.0
+ pdiblcb = -0.0001934
+ drout = 0.5264
+ pscbe1 = 5.12e+8
+ pscbe2 = 9.477e-8
+ pvag = 0.0
+ delta = 0.0457
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.016e-10
+ bgidl = 1.0e+9
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5162+sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_8}
+ kt2 = -0.122
+ at = 3.889e+4
+ ute = -0.3
+ ua1 = 1.346e-10
+ ub1 = 5.223e-19
+ uc1 = 6.005e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 10.0
+ xrcrg2 = 2.0
+ rbpb = {400*sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult}
+ rbpd = 0.001
+ rbps = 0.001
+ rbdb = 1.0e+5
+ rbsb = 1.0e+5
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = {1.25e-06+sky130_fd_pr__rf_pfet_01v8_b__xgw_diff}
+ xgl = 0.0
+ ngcon = 2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.363
+ jss = 2.148e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.002039
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.001241
+ tcjsw = 0.0003736
+ tcjswg = 0.001
+ cgdo = {1.3e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgso = {1e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.001e-11*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cgdl = {1.32e-10*sky130_fd_pr__rf_pfet_01v8_b__overlap_mult}
+ cf = 1.2e-11
+ clc = 0.0
+ cle = 0.6
+ dlc = {1e-09+sky130_fd_pr__rf_pfet_01v8_b__dlc_diff+sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__rf_pfet_01v8_b__dwc_diff}
+ vfbcv = -0.1447
+ acde = 0.401
+ moin = 15.0
+ noff = 2.5
+ voffcv = 0.05
+ ngate = 1.0e+23
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.002*sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult}
+ mjs = 0.1362
+ pbs = 0.9587
+ cjsws = {9.88e-11*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjsws = 0.92
+ pbsws = 0.94
+ cjswgs = {2.6e-10*sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult}
+ mjswgs = 0.12
+ pbswgs = 1.4
.ends sky130_fd_pr__rf_pfet_01v8_bM04W5p00
