* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 1
.param
+ sky130_fd_pr__special_pfet_01v8_hvt__toxe_mult = 0.9635
+ sky130_fd_pr__special_pfet_01v8_hvt__rshp_mult = 1.0
+ sky130_fd_pr__special_pfet_01v8_hvt__overlap_mult = 0.91216
+ sky130_fd_pr__special_pfet_01v8_hvt__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_pfet_01v8_hvt__wint_diff = -2.252e-8
+ sky130_fd_pr__special_pfet_01v8_hvt__dlc_diff = 1.21275e-8
+ sky130_fd_pr__special_pfet_01v8_hvt__dwc_diff = -2.252e-8
*
* sky130_fd_pr__special_pfet_01v8_hvt, Bin 000, W = 0.36, L = 0.15
* ------------------------------------
+ sky130_fd_pr__special_pfet_01v8_hvt__k2_diff_0 = -0.012919
+ sky130_fd_pr__special_pfet_01v8_hvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__ua_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__ub_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__ags_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__a0_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__voff_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__keta_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__b0_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__b1_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__vsat_diff_0 = 5500.8
+ sky130_fd_pr__special_pfet_01v8_hvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__u0_diff_0 = -0.00052794
+ sky130_fd_pr__special_pfet_01v8_hvt__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_01v8_hvt__vth0_diff_0 = 0.067192
*
.include "sky130_fd_pr__special_pfet_01v8_hvt__ff.pm3.spice"
