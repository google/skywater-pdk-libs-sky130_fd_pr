* Copyright 2022 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SKY130 Spice File.
.param
+ capunits = 1.0e-6
+ dkisepp5x = 0.745
+ dknfpp = 1.0
+ dknfpp5x = 1.0009
+ sky130_fd_pr__nfet_20v0_nvt_iso__k2_diff = -0.11937
+ sky130_fd_pr__nfet_20v0_nvt_iso__reverse_tmax = '20.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__reverse_vds = '-0.01'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbd_1 = '100.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbd_2 = '25.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbs_1 = '20.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_1 = '100.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_2 = '25.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgb_1 = '100.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgb_2 = '20.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgd_1 = 'sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgd_2 = 'sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_2'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgs_1 = '100.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgs_2 = '20.001n'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max_1 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max_2 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min_1 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min_2 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min - sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_reversemax = '0.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbd_reversemin = '-5.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max = '0.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max_1 = '0.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min = '-2.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1 = '-2.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_max = '22.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1 = '22.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2 = '22.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_min = '-0.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_min_1 = '-0.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vds_min_2 = '-0.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max_1 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1 - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max_2 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2 - sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min = '-1*sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max' + sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min_1 = '0 - 2.5'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min_2 = '0 - 2.5'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max_1 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max_2 = 'sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min = '-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min_1 = '-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min_2 = '-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemax = '5.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemax_1 = '0.101'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemin = '-5.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemin_1 = '-0.101'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max = '6.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1 = '5.751'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2 = '6.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min = '-1*6.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min_1 = '-1*5.751'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min_2 = '-1*6.001'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vsd_reversemax = '5.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vsd_reversemin = '-0.501'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vtx = '0.02'
+ sky130_fd_pr__special_nfet_pass_flash__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_pr__special_nfet_pass_flash__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__dwg_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt1l_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__lint_slope = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_slope = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nlx_diff = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__tox_slope = 0.006589
+ sky130_fd_pr__special_nfet_pass_flash__voff_slope = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__vth0_slope = 0.010889
+ sky130_fd_pr__special_nfet_pass_flash__wint_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_lint_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope = 0.12
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope = 0.008
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1 = 0.0205
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope2 = 0.01
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope3 = 0.0067
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope = 0.13
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_vth0_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__b_wint_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__lint1_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__lint_slope = 3.0e-9
+ sky130_fd_pr__rf_nfet_g5v0d10v5__nfactor_slope = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__tox2_slope = 0.0086
+ sky130_fd_pr__rf_nfet_g5v0d10v5__tox3_slope = 0.0055
+ sky130_fd_pr__rf_nfet_g5v0d10v5__tox4_slope = 0.0255
+ sky130_fd_pr__rf_nfet_g5v0d10v5__tox_offset = 0.0
+ sky130_fd_pr__rf_nfet_g5v0d10v5__tox_slope = 0.008
+ sky130_fd_pr__rf_nfet_g5v0d10v5__voff2_slope = 0.0085
+ sky130_fd_pr__rf_nfet_g5v0d10v5__voff_slope = 0.00375
+ sky130_fd_pr__rf_nfet_g5v0d10v5__wint_slope = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__b_toxe_slope = 0.003443
+ sky130_fd_pr__rf_nfet_01v8_lvt__b_vth0_slope = 0.006056
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__base__dlc_rotweak = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__toxe1_slope = 0.008089
+ sky130_fd_pr__rf_nfet_01v8_lvt__toxe_slope = 0.006789
+ sky130_fd_pr__special_nfet_pass_lvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_lvt__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_lvt__ua_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_lvt__ub_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_pass__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__kt1l_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__lint_slope = 0.0
+ sky130_fd_pr__special_nfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__nfactor_slope = 0.0
+ sky130_fd_pr__special_nfet_pass__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__tox_slope = 0.003589
+ sky130_fd_pr__special_nfet_pass__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__voff_slope = 0.0
+ sky130_fd_pr__special_nfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__vth0_slope = 0.005589
+ sky130_fd_pr__special_nfet_pass__wint_slope = 0.0
+ sky130_fd_pr__special_nfet_pass_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_latch__cdsc_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cdscb_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cdscd_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__cit_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_nfet_latch__dvt0_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__dvt1_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__kt2_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__lint_slope = 0.0
+ sky130_fd_pr__special_nfet_latch__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__nfactor_slope = 0.0
+ sky130_fd_pr__special_nfet_latch__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__tox_slope = 0.005989
+ sky130_fd_pr__special_nfet_latch__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__voff_slope = 0.0
+ sky130_fd_pr__special_nfet_latch__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__vth0_slope = 0.005289
+ sky130_fd_pr__special_nfet_latch__wint_slope = 0.0
+ sky130_fd_pr__special_nfet_latch_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__rf_nfet_01v8__b_toxe_slope = 0.003443
+ sky130_fd_pr__rf_nfet_01v8__b_voff_slope = 0.007
+ sky130_fd_pr__rf_nfet_01v8__b_vth0_slope = 0.005556
+ sky130_fd_pr__rf_nfet_01v8_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8__lint1_slope = 0.0
+ sky130_fd_pr__rf_nfet_01v8__lint_slope = 5.767e-9
+ sky130_fd_pr__rf_nfet_01v8__toxe1_slope = 0.006989
+ sky130_fd_pr__rf_nfet_01v8__toxe2_slope = 0.005989
+ sky130_fd_pr__rf_nfet_01v8__toxe3_slope = 0.01089
+ sky130_fd_pr__rf_nfet_01v8__toxe4_slope = 0.01289
+ sky130_fd_pr__rf_nfet_01v8__toxe_slope = 0.008989
+ sky130_fd_pr__special_pfet_pass__cdsc_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cdscb_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cdscd_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__cit_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__dlc_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__special_pfet_pass__dvt0_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__dwc_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__kt1l_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__kt2_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__lint_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__lint_slope = 0.0
+ sky130_fd_pr__special_pfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__nfactor_slope = 0.0
+ sky130_fd_pr__special_pfet_pass__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__tox_mult = 1.0
+ sky130_fd_pr__special_pfet_pass__tox_slope = 0.005567
+ sky130_fd_pr__special_pfet_pass__voff_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__voff_slope = 0.0
+ sky130_fd_pr__special_pfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__vth0_slope = 0.005567
+ sky130_fd_pr__special_pfet_pass__wint_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__wint_slope = 0.0
+ sky130_fd_pr__special_pfet_pass_lowleakage__dlc_rotweak = lv_dlc_rotweak
+ sky130_fd_pr__rf_pfet_01v8__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_pfet_01v8__aw_rs_mult = 1.0
+ sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1 = 0.1
+ sky130_fd_pr__rf_pfet_01v8__b_toxe_slope = 0.006443
+ sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1 = 0.004443
+ sky130_fd_pr__rf_pfet_01v8__b_voff_slope = 0.014
+ sky130_fd_pr__rf_pfet_01v8__b_voff_slope1 = 0.009
+ sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1 = 0.007356
+ sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2 = 0.009356
+ sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3 = 0.008356
+ sky130_fd_pr__rf_pfet_01v8_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8__nfactor1_slope = 0.0
+ sky130_fd_pr__rf_pfet_01v8__nfactor_slope = 0.429
+ sky130_fd_pr__rf_pfet_01v8__toxe1_slope = 0.01067
+ sky130_fd_pr__rf_pfet_01v8__toxe2_slope = 0.01167
+ sky130_fd_pr__rf_pfet_01v8__toxe3_slope = 0.01367
+ sky130_fd_pr__rf_pfet_01v8__toxe4_slope = 0.01467
+ sky130_fd_pr__rf_pfet_01v8__toxe5_slope = 0.01567
+ sky130_fd_pr__rf_pfet_01v8__toxe_slope = 0.01267
+ sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__dlc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_bs_flash__special_sonosfet_star__dwc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__k2_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0 = -0.44275
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_1 = -0.3267
+ sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_2 = -0.67944
+ sky130_fd_bs_flash__special_sonosfet_star__lint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__overlap_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__tox_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_star__tox_slope = 0.002
+ sky130_fd_bs_flash__special_sonosfet_star__tox_slope1 = 0.002
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0 = -0.0069221
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_1 = -0.0041919
+ sky130_fd_bs_flash__special_sonosfet_star__u0_diff_2 = -0.0081788
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__voff_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0 = 0.91203
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_1 = 1.3659
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_2 = 0.27494
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_slope = 0.0255
+ sky130_fd_bs_flash__special_sonosfet_star__vth0_slope1 = 0.028
+ sky130_fd_bs_flash__special_sonosfet_star__wint_diff = 0.0
+ sonos_eeol_dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_bs_flash__special_sonosfet_original__ajunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_original__dlc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__dlc_rotweak = hv_dlc_rotweak
+ sky130_fd_bs_flash__special_sonosfet_original__dwc_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__k2_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__k2_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__k2_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_0 = -0.36466
+ sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_1 = -0.029107
+ sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_2 = -0.65907
+ sky130_fd_bs_flash__special_sonosfet_original__lint_diff = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_0 = -0.23845
+ sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_1 = 1.3597
+ sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_2 = 1.0202
+ sky130_fd_bs_flash__special_sonosfet_original__overlap_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_original__pjunction_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__tox_mult = 1.0
+ sky130_fd_bs_flash__special_sonosfet_original__tox_slope = 0.005
+ sky130_fd_bs_flash__special_sonosfet_original__u0_diff_0 = -0.004
+ sky130_fd_bs_flash__special_sonosfet_original__u0_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__u0_diff_2 = 0.0013468
+ sky130_fd_bs_flash__special_sonosfet_original__voff_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__voff_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__voff_diff_2 = -0.20912
+ sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_0 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_1 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_2 = 0.0
+ sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_0 = -1.0278
+ sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_1 = -0.85561
+ sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_2 = -0.15565
+ sky130_fd_bs_flash__special_sonosfet_original__vth0_slope = 0.026
+ sky130_fd_bs_flash__special_sonosfet_original__wint_diff = 0.0
+ sonos_peol_dlc_rotweak = hv_dlc_rotweak
