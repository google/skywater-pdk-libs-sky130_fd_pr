* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 2
.param
+ sky130_fd_pr__special_nfet_01v8__toxe_mult = 0.948
+ sky130_fd_pr__special_nfet_01v8__rshn_mult = 1.0
+ sky130_fd_pr__special_nfet_01v8__overlap_mult = 0.94816
+ sky130_fd_pr__special_nfet_01v8__lint_diff = 1.21275e-8
+ sky130_fd_pr__special_nfet_01v8__wint_diff = -3.2175e-8
+ sky130_fd_pr__special_nfet_01v8__dlc_diff = 12.773e-9
+ sky130_fd_pr__special_nfet_01v8__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__special_nfet_01v8, Bin 000, W = 0.36, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_01v8__ub_diff_0 = 4.16095e-19
+ sky130_fd_pr__special_nfet_01v8__eta0_diff_0 = 3.2537e-5
+ sky130_fd_pr__special_nfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vsat_diff_0 = -65067.0
+ sky130_fd_pr__special_nfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vth0_diff_0 = -0.12224
+ sky130_fd_pr__special_nfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b0_diff_0 = -7.39989e-7
+ sky130_fd_pr__special_nfet_01v8__b1_diff_0 = 2.7011e-8
+ sky130_fd_pr__special_nfet_01v8__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pclm_diff_0 = 0.00091873
+ sky130_fd_pr__special_nfet_01v8__u0_diff_0 = -0.0083504
+ sky130_fd_pr__special_nfet_01v8__nfactor_diff_0 = 0.5935569
+ sky130_fd_pr__special_nfet_01v8__keta_diff_0 = 0.00306555
+ sky130_fd_pr__special_nfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_01v8__k2_diff_0 = 0.020341
+ sky130_fd_pr__special_nfet_01v8__ua_diff_0 = -4.02468e-11
*
* sky130_fd_pr__special_nfet_01v8, Bin 001, W = 0.39, L = 0.15
* -----------------------------------
+ sky130_fd_pr__special_nfet_01v8__ua_diff_1 = -4.99625e-12
+ sky130_fd_pr__special_nfet_01v8__ub_diff_1 = 3.05799e-19
+ sky130_fd_pr__special_nfet_01v8__eta0_diff_1 = 1.15988e-5
+ sky130_fd_pr__special_nfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vsat_diff_1 = -59191.0
+ sky130_fd_pr__special_nfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__vth0_diff_1 = -0.12953
+ sky130_fd_pr__special_nfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__b0_diff_1 = -4.77112e-7
+ sky130_fd_pr__special_nfet_01v8__b1_diff_1 = 2.47721e-8
+ sky130_fd_pr__special_nfet_01v8__voff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__pclm_diff_1 = 0.00032751
+ sky130_fd_pr__special_nfet_01v8__u0_diff_1 = -0.0072906
+ sky130_fd_pr__special_nfet_01v8__nfactor_diff_1 = 0.56383409
+ sky130_fd_pr__special_nfet_01v8__keta_diff_1 = 0.0010928
+ sky130_fd_pr__special_nfet_01v8__ags_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_01v8__k2_diff_1 = 0.022274
*
.include "sky130_fd_pr__special_nfet_01v8__sf.pm3.spice"
