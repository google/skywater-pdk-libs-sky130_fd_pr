* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
* 	mismatch {
*     	}
* }
.subckt  sky130_fd_pr__res_high_po_5p73 r0 r1 b
+ 
.param  w = 5.730 l = 5 mult = 1.0
+ 
+ body_pelgrom = 0.037
+ rend_mm = 0.01
+ rcon = 68.05
+ rsheet = 56.46
+ tc1_voltco = 2.35e-2
+ vc1_body = -2.62e-5
+ vc2_body = 2.25e-5
+ vc1_raw_end = 8.74e-4
+ vc2_raw_end = -1.34e-2
+ vc3_raw_end = 1.72e-2
+ r0_var = 4.29
+ r1_var = 1.6
+ vc1_end = {vc1_raw_end*2.865/l*(1+(tc1_voltco*min((temp-30),0)))}
+ vc2_end = {vc2_raw_end*2.865/l*(1+(tc1_voltco*min((temp-30),0)))}
+ vc3_end = {vc3_raw_end*2.865/l*(1+(tc1_voltco*min((temp-30),0)))}
+ rtot_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2*pow(r0_var,2)+pow((r1_var*l),2))}
+ rend_var = {sky130_fd_pr__res_high_po__var_mult*sqrt(2)*r0_var}
+ rbody_var = {rtot_var-rend_var}
+ res_match = {(body_pelgrom/sqrt(w*l*mult))*sky130_fd_pr__res_high_po__slope_spectre}
+ rend = {(rcon+rend_var)*(1+rend_mm/sqrt(mult)*sky130_fd_pr__res_high_po__con_slope_spectre)}
+ rbody = {(l*rsheet+rbody_var)*(1+res_match)}
rend r0 ra r = {rend*(1+min(abs(v(r0,r1)),2.0)*vc1_end+pow(min(abs(v(r0,r1)),2.0),2)*vc2_end+pow(min(abs(v(r0,r1)),2.0),3)*vc3_end)}
rhrpoly_5p73 ra r1 resbody r = {rbody*(1+abs(v(r0,r1))*vc1_body+pow(abs(v(r0,r1)),2)*vc2_body)}
c1 r0 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_16_2*1e-6)/2}
c2 r1 b c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_16_2*1e-6)/2}
.model resbody r tc1 = {tc1rpolybody} tc2 = {tc2rpolybody} tnom = 30.0
.ends sky130_fd_pr__res_high_po_5p73
