* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_nfet_pass_lvt__tox_slope_spectre = 0.0
.param sky130_fd_pr__special_nfet_pass_lvt__vth0_slope_spectre = 0.0
* statistics {
*   mismatch {
*     vary sky130_fd_pr__special_nfet_pass_lvt__tox_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_pass_lvt__vth0_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__special_nfet_pass_lvt d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 mult = 1 sa = 0 sb = 0 sd = 0.0
msky130_fd_pr__special_nfet_pass_lvt d g s b sky130_fd_pr__special_nfet_pass_lvt__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs}
.model sky130_fd_pr__special_nfet_pass_lvt__model.0 nmos
* Model Flag Parameters
+ lmin = 1.45e-007 lmax = 1.55e-007 wmin = 2.95e-007 wmax = 3.05e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__special_nfet_pass_lvt__tox_slope_spectre)
+ toxe = {4.148e-009*sky130_fd_pr__special_nfet_pass_lvt__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*4.148e-09*2.443e-3*sky130_fd_pr__special_nfet_pass_lvt__toxe_mult/sqrt(l*w*mult)}
+ toxm = 4.148e-9
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1*sky130_fd_pr__special_nfet_pass_lvt__rshn_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {2.6e-008+sky130_fd_pr__special_nfet_pass_lvt__wint_diff}
+ lint = {1.2025e-008+sky130_fd_pr__special_nfet_pass_lvt__lint_diff}
*(mismatch parameter sky130_fd_pr__special_nfet_pass_lvt__vth0_slope_spectre)
+ vth0 = {0.41207609+sky130_fd_pr__special_nfet_pass_lvt__vth0_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*5.456e-03/sqrt(l*w*mult)}
+ k1 = 0.5273401
+ k2 = {-0.019324124+sky130_fd_pr__special_nfet_pass_lvt__k2_diff_0}
+ k3 = 1.65
+ k3b = 1.6
+ w0 = 1.0e-7
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ dsub = 0.24915505
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = -0.2
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 1.5e-5
+ cit = 9.9e-8
+ voff = {-0.15+sky130_fd_pr__special_nfet_pass_lvt__voff_diff_0}
+ nfactor = {1.7244198+sky130_fd_pr__special_nfet_pass_lvt__nfactor_diff_0}
+ eta0 = {0.067583862+sky130_fd_pr__special_nfet_pass_lvt__eta0_diff_0}
+ etab = -0.013910732
+ vfb = 0.0
+ u0 = {0.046750961+sky130_fd_pr__special_nfet_pass_lvt__u0_diff_0}
+ ua = {5e-11+sky130_fd_pr__special_nfet_pass_lvt__ua_diff_0}
+ ub = {4e-19+sky130_fd_pr__special_nfet_pass_lvt__ub_diff_0}
+ uc = -2.7110648e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 0.0
+ vsat = {151538.73+sky130_fd_pr__special_nfet_pass_lvt__vsat_diff_0}
+ a0 = 1.0
+ ags = 15.0
+ a1 = 0.0
+ a2 = 0.38689047
+ b0 = 0.0
+ b1 = 0.0
+ keta = 0.05
+ dwg = -1.33e-8
+ dwb = -1.08e-8
+ pclm = 0.47255423
+ pdiblc1 = 9.9e-13
+ pdiblc2 = 9.9e-13
+ pdiblcb = -0.1
+ drout = 0.9999
+ pscbe1 = 8.0476145e+8
+ pscbe2 = 9.9022619e-9
+ pvag = 0.0018113134
+ delta = 0.01
+ fprout = 3.289058e-11
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 168.29597
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 9.9e-6
+ prwg = 0.0
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.01
+ alpha1 = 1.9991339
+ beta0 = 33.32325
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
* Charge AND Capacitance Model Parameters
+ dlc = {1.3469e-008+sky130_fd_pr__special_nfet_pass_lvt__dlc_diff}
+ dwc = {2.6e-008+sky130_fd_pr__special_nfet_pass_lvt__dwc_diff}
+ xpart = 0.0
+ cgso = {2.5889e-010*sky130_fd_pr__special_nfet_pass_lvt__overlap_mult}
+ cgdo = {2.5889e-010*sky130_fd_pr__special_nfet_pass_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ cgdl = {2.5e-011*sky130_fd_pr__special_nfet_pass_lvt__overlap_mult}
+ cgsl = {2.5e-011*sky130_fd_pr__special_nfet_pass_lvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.0e-14
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
* High-Speed/RF Model Parameters
* Flicker AND Thermal Noise Model Parameters
+ ef = 1.2
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 8.0e+11
+ em = 4.1e+7
+ lintnoi = -3.0e-7
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
+ rnoia = 0.912
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.9
+ xjbvs = 1.0
+ pbs = 0.7477
+ cjs = {0.001209*sky130_fd_pr__special_nfet_pass_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbsws = 0.1
+ cjsws = {3.6224e-011*sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbswgs = 0.79644
+ cjswgs = {2.0132e-010*sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult}
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.18424344
+ kt2 = -0.021488214
+ at = 33001.301
+ ute = -1.7796658
+ ua1 = -1.914008e-10
+ ub1 = 3.9161781e-19
+ uc1 = 1.8902599e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.195e-6
+ sbref = 2.585e-6
+ kvth0 = 7.9e-9
+ lkvth0 = 0.0
+ wkvth0 = 3.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.ends sky130_fd_pr__special_nfet_pass_lvt
