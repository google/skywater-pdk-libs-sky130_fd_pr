* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./models_global.spice created from ./models.spice
*
***********************************
* Model dimensions are in um:
* ---------------------------------

.option scale=1.0u
.options parser scale=1.0u


***********************************
* Global parameter values
* ---------------------------------

.param
+ sw_tox_lv_nom = 4.148E-09
+ sw_tox_hv_nom = 11.60E-09


***********************************
* Global functions
* ---------------------------------

.param
* Separate Tox Corners from Monte Carlo for fet ff and ss
+ sw_tox_lv = {sw_tox_lv_corner+sw_tox_lv_mc}
+ sw_tox_hv = {sw_tox_hv_corner+sw_tox_hv_mc}
+ sw_func_tox_lv_ratio = {sw_tox_lv/sw_tox_lv_nom}
+ sw_func_tox_hv_ratio = {sw_tox_hv/sw_tox_hv_nom}
+ sw_func_nsd_pw_cj = {sw_nsd_pw_cj/1.35E-03}
+ sw_func_psd_nw_cj = {sw_psd_nw_cj/7.3802e-4}
+ sw_func_nw_pw_cj = {sw_nw_pw_cj/9.000e-5}
+ sw_func_pw_dnw_cj = {sw_pw_dnw_cj/3.824e-4}
+ sw_func_dnw_sub_cj = {sw_dnw_sub_cj/7.743e-5}
+ sw_func_rdp = {sw_rdp/197}
+ sw_func_rdn = {sw_rdn/120}
+ sw_func_pw_rs = {sw_pw_rs/3816}


*************************************************************
* Matching constants.
*    Note: Between two device mismatch:
*	                                Matching Constant * sqrt(2/dimension)
* -----------------------------------------------------------

.param
+ sw_mm_tox_lv = {3.443e-03*sw_tox_lv_nom} ;  41A  gate oxide 
+ sw_mm_tox_hv = {5.800e-03*sw_tox_hv_nom} ;  116A gate oxide
+ sw_mm_vth0_sky130_fd_pr__nfet_01v8 = 3.356e-03 ;  Nmos VT
+ sw_mm_vth0_sky130_fd_pr__nfet_01v8_lvt = 5.456e-03 ;  Nmos LowVt VT
+ sw_mm_vth0_sky130_fd_pr__nfet_g5v0d10v5 = 8.200e-03 ;  5V Nmos VT, data 11.6/sqrt(2)
+ sw_mm_vth0_sky130_fd_pr__nfet_01v8_nat = 6.000e-03 ;  Native VT, was 1.2e-3 seemed too low
+ sw_mm_vth0_sky130_fd_pr__nfet_g5v0d16v0 = 8.000e-03 ;  12V Nmos VT, original was 0.8, too high
+ sw_mm_vth0_sky130_fd_pr__pfet_01v8 = 5.856e-03 ;  Pmos VT
+ sw_mm_vth0_sky130_fd_pr__pfet_01v8_lvt = 1.089e-02 ;  Pmos LowVt VT
+ sw_mm_vth0_sky130_fd_pr__pfet_01v8_hvt = 5.500e-03 ;  Pmos HighVt VT
+ sw_mm_vth0_sky130_fd_pr__pfet_g5v0d10v5 = 1.200e-02 ;  5V Pmos VT, estimated, was zero
+ sw_mm_vth0_sky130_fd_pr__pfet_g5v0d16v0 = 1.200e-02 ;  12V Pmos VT, was 0.0 
+ sw_mm_cmim = 4.700e-03 ;  MIM capacitor Ca CBCM data
+ sw_mm_cvpp = 9.000e-03 ;  Vertical Plate capacitors
+ sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_bf = 5.537e-02 ;  PNP BF
+ sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_is = 1.662e-02 ;  PNP IS
+ sw_mm_npn_bf = 5.000e-02 ;  NPN BF
+ sw_mm_npn_is = 3.000e-03 ;  NPN IS
+ sw_mm_sky130_fd_pr__res_iso_pw = 1.000e-02 ;  Pwell resistor, estimated
+ sw_mm_sky130_fd_pr__res_generic_po = 1.200e-01 ;  50 Ohm-sq Poly resistor
+ sw_mm_sky130_fd_pr__res_high_po = 2.060e-02 ;  300 Ohm-sq Poly resistor (data), was 3.552e-2 (Cypress)
+ sw_mm_sky130_fd_pr__res_xhigh_po = 4.640e-02 ;  2K  Ohm-sq Poly resistor (based on data)
+ sw_mm_sky130_fd_pr__res_generic_po_head = 6.300e-02 ;  Poly resistor head


************************************
* Global Matching Monte Carlo driver
* ----------------------------------

.param mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1) = 0 mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1) = 0
*    statistics{
*       mismatch{
*          vary mm_z1 dist=gauss std=mismatch_factor
*          vary mm_z2 dist=gauss std=mismatch_factor
*       }
*    }


************************************
* Process Monte Carlo
*    Log Normal std = ln(std ratio)*ln(mean)
* ----------------------------------

*  Independent arameters used to Monte Carlo only (*_mc)
*  The remaining parameters are used both Corners and MC.
.param
+ sw_tox_lv_mc = 0
+ sw_tox_hv_mc = 0
+ sw_vth0_sky130_fd_pr__nfet_01v8_lvt_mc = 0
+ sw_pw_rs_mc = 1
+ sw_vth0_sky130_fd_pr__nfet_01v8_mc = 0
+ sw_vth0_sky130_fd_pr__pfet_01v8_lvt_mc = 0
+ sw_vth0_sky130_fd_pr__pfet_01v8_hvt_mc = 0
+ sw_vth0_sky130_fd_pr__pfet_01v8_mc = 0
+ sw_vth0_sky130_fd_pr__nfet_01v8_nat_mc = 0
+ sw_vth0_sky130_fd_pr__nfet_g5v0d10v5_mc = 0
+ sw_vth0_sky130_fd_pr__pfet_g5v0d10v5_mc = 0
+ sw_vth0_sky130_fd_pr__nfet_g5v0d16v0_mc = 0
+ sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc = 0
*  ----------------------------


*    statistics{
*       process{
*          vary sw_tox_lv_mc             dist=gauss   std=0.375e-10*process_mc_factor
*          vary sw_tox_hv_mc             dist=gauss   std=1.25e-10*process_mc_factor
*          vary sw_polycd                dist=gauss   std=1.5e-9*process_mc_factor
*          vary sw_activecd              dist=gauss   std=5.0e-9*process_mc_factor
*          vary sw_fox_cap               dist=gauss   std=0.0475*process_mc_factor
*          vary sw_li_cap                dist=lnorm   std=0.1*process_mc_factor
*          vary sw_fox_poly_cap          dist=gauss   std=0.0475*process_mc_factor
*          vary sw_nw_rs_mult            dist=lnorm   std=0.12*process_mc_factor
*          vary sw_pw_rs_mc              dist=gauss   std=6.6*process_mc_factor       percent=yes
*          vary sw_nldd                  dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_nsd_pw_cj             dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_psd_nw_cj             dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_nw_pw_cj              dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_pw_dnw_cj             dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_dnw_sub_cj            dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_vth0_sky130_fd_pr__nfet_01v8_mc          dist=gauss   std=0.006*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__nfet_01v8_lvt_mc      dist=gauss   std=0.006*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__nfet_g5v0d10v5_mc       dist=gauss   std=0.010*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__nfet_01v8_nat_mc      dist=gauss   std=0.006*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__nfet_g5v0d16v0_mc   dist=gauss   std=0.035*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__nfet_01v8_zvt         dist=gauss   std=0.007*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__pfet_01v8_mc          dist=gauss   std=0.009*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__pfet_01v8_lvt_mc      dist=gauss   std=0.023*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__pfet_01v8_hvt_mc      dist=gauss   std=0.009*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__pfet_g5v0d10v5_mc       dist=gauss   std=0.02*process_mc_factor
*          vary sw_vth0_sky130_fd_pr__pfet_g5v0d16v0_mc   dist=gauss   std=0.03*process_mc_factor
*          vary sw_cap_mim_ca            dist=gauss   std=2.7*process_mc_factor       percent=yes
*          vary sw_cap_mim_dw            dist=gauss   std=24e-9*process_mc_factor
*          vary sw_sky130_fd_pr__res_generic_m1_rs                dist=gauss   std=5*process_mc_factor         percent=yes
*          vary sw_sky130_fd_pr__res_generic_m2_rs                dist=gauss   std=5*process_mc_factor         percent=yes
*          vary sw_sky130_fd_pr__res_generic_m3_rs                dist=gauss   std=5*process_mc_factor         percent=yes
*          vary sw_sky130_fd_pr__res_generic_m4_rs                dist=gauss   std=5*process_mc_factor         percent=yes
*          vary sw_m3_dw                 dist=gauss   std=1.6e-8*process_mc_factor
*          vary sw_m4_dw                 dist=gauss   std=1.6e-8*process_mc_factor
*          vary sw_rcvia                 dist=lnorm   std=0.26*process_mc_factor
*          vary sw_rcvia2                dist=lnorm   std=0.21*process_mc_factor
*          vary sw_rcvia3                dist=lnorm   std=0.21*process_mc_factor
*          vary sw_rcvia4                dist=lnorm   std=0.21*process_mc_factor
*          vary sw_rcl1                  dist=lnorm   std=0.39*process_mc_factor
*          vary sw_rl1                   dist=gauss   std=5*process_mc_factor         percent=yes
*          vary sw_rnw                   dist=gauss   std=3.75*process_mc_factor      percent=yes 
*          vary sw_rp1                   dist=gauss   std=2.5*process_mc_factor       percent=yes 
*          vary sw_rcn                   dist=lnorm   std=0.9*process_mc_factor         
*          vary sw_rcp1                  dist=lnorm   std=0.86*process_mc_factor
*          vary sw_rdp                   dist=gauss   std=3.75*process_mc_factor      percent=yes
*          vary sw_rdn                   dist=gauss   std=2.5*process_mc_factor       percent=yes
*          vary sw_poly_head_res         dist=gauss   std=2.5*process_mc_factor       percent=yes 
*          vary sw_sky130_fd_pr__res_high_po_rs           dist=gauss   std=3.5*process_mc_factor       percent=yes
*          vary sw_sky130_fd_pr__res_xhigh_po_rs         dist=gauss   std=4.0*process_mc_factor       percent=yes     
*       }
*    }


********************************************************
********End of global parameters and definitions *******
********************************************************
********************************************************
********************************************************



