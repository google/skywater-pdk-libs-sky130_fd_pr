* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./parameters_res_high.spice created from ./parameters.spice
*
.param sw_sky130_fd_pr__res_high_po_rs = {325.0+corner_factor*45.0} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.035,1)
.param sw_sky130_fd_pr__res_xhigh_po_rs = {2000.0+corner_factor*300.0} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.04,1)
.param sw_poly_head_res = {1.0+corner_factor*0.125} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_sky130_fd_pr__res_generic_m1_rs = {0.124+corner_factor*0.01899999999999999} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.05,1)
.param sw_sky130_fd_pr__res_generic_m2_rs = {0.124+corner_factor*0.01899999999999999} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.05,1)
.param sw_sky130_fd_pr__res_generic_m3_rs = {0.046+corner_factor*0.006999999999999999} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.05,1)
.param sw_sky130_fd_pr__res_generic_m4_rs = {0.046+corner_factor*0.006999999999999999} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.05,1)
.param sw_sky130_fd_pr__res_generic_m5_rs = {0.0275+corner_factor*0.0045000000000000005}
.param sw_m1_dw = {0.0+corner_factor*-2.5e-08}
.param sw_m2_dw = {0.0+corner_factor*-2.5e-08}
.param sw_m3_dw = {0.0+corner_factor*-6.5e-08} + process_mc_factor*MC_PR_SWITCH*AGAUSS(0,1.6e-08,1)
.param sw_m4_dw = {0.0+corner_factor*-6.5e-08} + process_mc_factor*MC_PR_SWITCH*AGAUSS(0,1.6e-08,1)
.param sw_m5_dw = {0.0+corner_factor*-1.7e-07}
.param sw_rcvia = {4.5+corner_factor*7.35} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.26,1))
.param sw_rcvia2 = {3.41+corner_factor*3.213} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.21,1))
.param sw_rcvia3 = {3.41+corner_factor*3.213} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.21,1))
.param sw_rcvia4 = {3.41+corner_factor*3.213} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.21,1))
.param sw_rcl1 = {9.3+corner_factor*9.309999999999999} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.39,1))
.param sw_rl1 = {12.3+corner_factor*2.5} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.05,1)
.param sw_rl1_dw = {0.0+corner_factor*-2e-08}
.param sw_rnw = {1700.0+corner_factor*460.0} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.0375,1)
.param sw_rp1 = {48.2+corner_factor*7.399999999999999} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_rcn = {182.0+corner_factor*114.0} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.9,1))
.param sw_rcp1 = {145.0+corner_factor*84.0} + process_mc_factor*MC_PR_SWITCH*EXP(AGAUSS(0,0.86,1))
.param sw_rdn = {120.0+corner_factor*12.0} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.025,1)
.param sw_rdp = {197.0+corner_factor*31.0} + process_mc_factor*MC_PR_SWITCH*GAUSS(0,0.0375,1)
.param sw_pw_rs = {3816.0+corner_factor*1034.0}
