# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__fuse_m4__example1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__fuse_m4__example1 ;
  ORIGIN  0.800000  0.000000 ;
  SIZE  8.800000 BY  0.800000 ;
  OBS
    LAYER met3 ;
      RECT -0.800000 0.000000 0.000000 0.800000 ;
      RECT  7.200000 0.000000 8.000000 0.800000 ;
    LAYER met4 ;
      RECT -0.800000 0.000000 8.000000 0.800000 ;
    LAYER via3 ;
      RECT -0.560000 0.240000 -0.240000 0.560000 ;
      RECT  7.440000 0.240000  7.760000 0.560000 ;
  END
END sky130_fd_pr__fuse_m4__example1
END LIBRARY
