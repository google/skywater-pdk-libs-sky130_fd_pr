* SKY130 Spice File.
.include "all.spice"
.include "ff/legacy.spice"
.include "ff/nonfet.spice"
.include "ff/rf.spice"
