# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__padplhp__example_179573804
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__padplhp__example_179573804 ;
  ORIGIN  2.700000  2.700000 ;
  SIZE  65.40000 BY  65.40000 ;
  OBS
    LAYER met4 ;
      POLYGON -2.700000  3.830000 -2.280000  3.830000 -2.280000  3.410000 ;
      POLYGON -2.690000 56.180000 -2.690000 56.170000 -2.700000 56.170000 ;
      POLYGON -2.645000 56.225000 -2.645000 56.180000 -2.690000 56.180000 ;
      POLYGON -2.280000  3.410000 -1.100000  3.410000 -1.100000  2.230000 ;
      POLYGON -1.100000  2.230000 -0.680000  2.230000 -0.680000  1.810000 ;
      POLYGON -1.030000 57.840000 -1.030000 56.225000 -2.645000 56.225000 ;
      POLYGON -0.680000  1.810000  0.500000  1.810000  0.500000  0.630000 ;
      POLYGON  0.000000  4.950000  1.540000  3.410000  0.000000  3.410000 ;
      POLYGON  0.000000 56.180000  1.130000 56.180000  0.000000 55.050000 ;
      POLYGON  0.500000  0.630000  1.130000  0.630000  1.130000  0.000000 ;
      POLYGON  0.570000 59.440000  0.570000 57.840000 -1.030000 57.840000 ;
      POLYGON  1.130000  0.000000  2.100000  0.000000  2.100000 -0.970000 ;
      POLYGON  1.130000 58.260000  3.210000 58.260000  1.130000 56.180000 ;
      POLYGON  1.130000 60.000000  1.130000 59.440000  0.570000 59.440000 ;
      POLYGON  1.540000  3.410000  3.140000  1.810000  1.540000  1.810000 ;
      POLYGON  2.100000 -0.970000  2.530000 -0.970000  2.530000 -1.400000 ;
      POLYGON  2.170000 61.040000  2.170000 60.000000  1.130000 60.000000 ;
      POLYGON  2.530000 -1.400000  3.710000 -1.400000  3.710000 -2.580000 ;
      POLYGON  3.140000  1.810000  3.820000  1.130000  3.140000  1.130000 ;
      POLYGON  3.210000 59.440000  4.390000 59.440000  3.210000 58.260000 ;
      POLYGON  3.710000 -2.580000  3.830000 -2.580000  3.830000 -2.700000 ;
      POLYGON  3.820000  1.130000  4.950000  0.000000  3.820000  0.000000 ;
      POLYGON  3.830000 62.700000  3.830000 61.040000  2.170000 61.040000 ;
      POLYGON  4.390000 59.860000  4.810000 59.860000  4.390000 59.440000 ;
      POLYGON  4.810000 60.000000  4.950000 60.000000  4.810000 59.860000 ;
      POLYGON 55.050000 60.000000 55.190000 60.000000 55.190000 59.860000 ;
      POLYGON 55.190000 59.860000 55.260000 59.860000 55.260000 59.790000 ;
      POLYGON 55.260000 59.790000 55.610000 59.790000 55.610000 59.440000 ;
      POLYGON 55.610000 59.440000 55.680000 59.440000 55.680000 59.370000 ;
      POLYGON 55.680000 59.370000 56.790000 59.370000 56.790000 58.260000 ;
      POLYGON 56.170000 -1.040000 57.830000 -1.040000 56.170000 -2.700000 ;
      POLYGON 56.170000 62.700000 56.290000 62.580000 56.170000 62.580000 ;
      POLYGON 56.180000  1.130000 56.180000  0.000000 55.050000  0.000000 ;
      POLYGON 56.290000 62.580000 57.900000 60.970000 56.290000 60.970000 ;
      POLYGON 56.790000  1.740000 56.790000  1.130000 56.180000  1.130000 ;
      POLYGON 56.790000 58.260000 56.860000 58.260000 56.860000 58.190000 ;
      POLYGON 56.860000  1.810000 56.860000  1.740000 56.790000  1.740000 ;
      POLYGON 56.860000 58.190000 57.280000 58.190000 57.280000 57.770000 ;
      POLYGON 57.280000 57.770000 58.460000 57.770000 58.460000 56.590000 ;
      POLYGON 57.830000  0.000000 58.870000  0.000000 57.830000 -1.040000 ;
      POLYGON 57.900000 60.970000 58.870000 60.000000 57.900000 60.000000 ;
      POLYGON 58.390000  3.340000 58.390000  1.810000 56.860000  1.810000 ;
      POLYGON 58.460000  3.410000 58.460000  3.340000 58.390000  3.340000 ;
      POLYGON 58.460000 56.590000 58.870000 56.590000 58.870000 56.180000 ;
      POLYGON 58.870000  0.560000 59.430000  0.560000 58.870000  0.000000 ;
      POLYGON 58.870000 56.180000 60.000000 56.180000 60.000000 55.050000 ;
      POLYGON 58.870000 60.000000 59.500000 59.370000 58.870000 59.370000 ;
      POLYGON 59.430000  1.740000 60.610000  1.740000 59.430000  0.560000 ;
      POLYGON 59.500000 59.370000 60.000000 58.870000 59.500000 58.870000 ;
      POLYGON 60.000000  4.950000 60.000000  3.410000 58.460000  3.410000 ;
      POLYGON 60.000000 58.870000 61.100000 57.770000 60.000000 57.770000 ;
      POLYGON 60.610000  2.160000 61.030000  2.160000 60.610000  1.740000 ;
      POLYGON 61.030000  3.340000 62.210000  3.340000 61.030000  2.160000 ;
      POLYGON 61.100000 57.770000 62.700000 56.170000 61.100000 56.170000 ;
      POLYGON 62.210000  3.775000 62.645000  3.775000 62.210000  3.340000 ;
      POLYGON 62.645000  3.830000 62.700000  3.830000 62.645000  3.775000 ;
      RECT -2.700000  3.830000  0.000000 56.170000 ;
      RECT -2.690000 56.170000  0.000000 56.180000 ;
      RECT -2.645000 56.180000  1.130000 56.225000 ;
      RECT -2.280000  3.410000  0.000000  3.830000 ;
      RECT -1.100000  2.230000  1.540000  3.410000 ;
      RECT -1.030000 56.225000  1.130000 57.840000 ;
      RECT -0.680000  1.810000  1.540000  2.230000 ;
      RECT  0.500000  0.630000  3.820000  1.130000 ;
      RECT  0.500000  1.130000  3.140000  1.810000 ;
      RECT  0.570000 57.840000  1.130000 58.260000 ;
      RECT  0.570000 58.260000  3.210000 59.440000 ;
      RECT  1.130000  0.000000  3.820000  0.630000 ;
      RECT  1.130000 59.440000  4.390000 59.860000 ;
      RECT  1.130000 59.860000  4.810000 60.000000 ;
      RECT  2.100000 -0.970000 57.830000  0.000000 ;
      RECT  2.170000 60.000000 57.900000 60.970000 ;
      RECT  2.170000 60.970000 56.290000 61.040000 ;
      RECT  2.530000 -1.400000 56.170000 -1.040000 ;
      RECT  2.530000 -1.040000 57.830000 -0.970000 ;
      RECT  3.710000 -2.580000 56.170000 -1.400000 ;
      RECT  3.830000 -2.700000 56.170000 -2.580000 ;
      RECT  3.830000 61.040000 56.290000 62.580000 ;
      RECT  3.830000 62.580000 56.170000 62.700000 ;
      RECT 55.190000 59.860000 58.870000 60.000000 ;
      RECT 55.260000 59.790000 58.870000 59.860000 ;
      RECT 55.610000 59.440000 58.870000 59.790000 ;
      RECT 55.680000 59.370000 58.870000 59.440000 ;
      RECT 56.180000  0.000000 58.870000  0.560000 ;
      RECT 56.180000  0.560000 59.430000  1.130000 ;
      RECT 56.790000  1.130000 59.430000  1.740000 ;
      RECT 56.790000 58.260000 60.000000 58.870000 ;
      RECT 56.790000 58.870000 59.500000 59.370000 ;
      RECT 56.860000  1.740000 60.610000  1.810000 ;
      RECT 56.860000 58.190000 60.000000 58.260000 ;
      RECT 57.280000 57.770000 60.000000 58.190000 ;
      RECT 58.390000  1.810000 60.610000  2.160000 ;
      RECT 58.390000  2.160000 61.030000  3.340000 ;
      RECT 58.460000  3.340000 62.210000  3.410000 ;
      RECT 58.460000 56.590000 61.100000 57.770000 ;
      RECT 58.870000 56.180000 61.100000 56.590000 ;
      RECT 60.000000  3.410000 62.210000  3.775000 ;
      RECT 60.000000  3.775000 62.645000  3.830000 ;
      RECT 60.000000  3.830000 62.700000 56.170000 ;
      RECT 60.000000 56.170000 61.100000 56.180000 ;
    LAYER met5 ;
      POLYGON -2.700000  3.830000 -2.280000  3.830000 -2.280000  3.410000 ;
      POLYGON -2.645000 56.225000 -2.645000 56.170000 -2.700000 56.170000 ;
      POLYGON -2.280000  3.410000 -1.100000  3.410000 -1.100000  2.230000 ;
      POLYGON -1.100000  2.230000 -0.680000  2.230000 -0.680000  1.810000 ;
      POLYGON -1.030000 57.840000 -1.030000 56.225000 -2.645000 56.225000 ;
      POLYGON -0.680000  1.810000  0.500000  1.810000  0.500000  0.630000 ;
      POLYGON  0.500000  0.630000  0.920000  0.630000  0.920000  0.210000 ;
      POLYGON  0.570000 59.440000  0.570000 57.840000 -1.030000 57.840000 ;
      POLYGON  0.920000  0.210000  2.100000  0.210000  2.100000 -0.970000 ;
      POLYGON  2.100000 -0.970000  2.530000 -0.970000  2.530000 -1.400000 ;
      POLYGON  2.170000 61.040000  2.170000 59.440000  0.570000 59.440000 ;
      POLYGON  2.530000 -1.400000  3.710000 -1.400000  3.710000 -2.580000 ;
      POLYGON  3.710000 -2.580000  3.830000 -2.580000  3.830000 -2.700000 ;
      POLYGON  3.830000 62.700000  3.830000 61.040000  2.170000 61.040000 ;
      POLYGON 56.170000 -1.040000 57.830000 -1.040000 56.170000 -2.700000 ;
      POLYGON 56.170000 62.700000 56.290000 62.580000 56.170000 62.580000 ;
      POLYGON 56.290000 62.580000 57.900000 60.970000 56.290000 60.970000 ;
      POLYGON 57.830000  0.140000 59.010000  0.140000 57.830000 -1.040000 ;
      POLYGON 57.900000 60.970000 59.500000 59.370000 57.900000 59.370000 ;
      POLYGON 59.010000  0.560000 59.430000  0.560000 59.010000  0.140000 ;
      POLYGON 59.430000  1.740000 60.610000  1.740000 59.430000  0.560000 ;
      POLYGON 59.500000 59.370000 61.100000 57.770000 59.500000 57.770000 ;
      POLYGON 60.610000  2.160000 61.030000  2.160000 60.610000  1.740000 ;
      POLYGON 61.030000  3.340000 62.210000  3.340000 61.030000  2.160000 ;
      POLYGON 61.100000 57.770000 62.700000 56.170000 61.100000 56.170000 ;
      POLYGON 62.210000  3.775000 62.645000  3.775000 62.210000  3.340000 ;
      POLYGON 62.645000  3.830000 62.700000  3.830000 62.645000  3.775000 ;
      RECT -2.700000  3.830000 62.700000 56.170000 ;
      RECT -2.645000 56.170000 61.100000 56.225000 ;
      RECT -2.280000  3.410000 62.210000  3.775000 ;
      RECT -2.280000  3.775000 62.645000  3.830000 ;
      RECT -1.100000  2.230000 61.030000  3.340000 ;
      RECT -1.100000  3.340000 62.210000  3.410000 ;
      RECT -1.030000 56.225000 61.100000 57.770000 ;
      RECT -1.030000 57.770000 59.500000 57.840000 ;
      RECT -0.680000  1.810000 60.610000  2.160000 ;
      RECT -0.680000  2.160000 61.030000  2.230000 ;
      RECT  0.500000  0.630000 59.430000  1.740000 ;
      RECT  0.500000  1.740000 60.610000  1.810000 ;
      RECT  0.570000 57.840000 59.500000 59.370000 ;
      RECT  0.570000 59.370000 57.900000 59.440000 ;
      RECT  0.920000  0.210000 59.010000  0.560000 ;
      RECT  0.920000  0.560000 59.430000  0.630000 ;
      RECT  2.100000 -0.970000 57.830000  0.140000 ;
      RECT  2.100000  0.140000 59.010000  0.210000 ;
      RECT  2.170000 59.440000 57.900000 60.970000 ;
      RECT  2.170000 60.970000 56.290000 61.040000 ;
      RECT  2.530000 -1.400000 56.170000 -1.040000 ;
      RECT  2.530000 -1.040000 57.830000 -0.970000 ;
      RECT  3.710000 -2.580000 56.170000 -1.400000 ;
      RECT  3.830000 -2.700000 56.170000 -2.580000 ;
      RECT  3.830000 61.040000 56.290000 62.580000 ;
      RECT  3.830000 62.580000 56.170000 62.700000 ;
    LAYER via4 ;
      RECT -2.580000  3.845000 -1.400000  5.025000 ;
      RECT -2.580000  5.445000 -1.400000  6.625000 ;
      RECT -2.580000  7.045000 -1.400000  8.225000 ;
      RECT -2.580000  8.645000 -1.400000  9.825000 ;
      RECT -2.580000 10.245000 -1.400000 11.425000 ;
      RECT -2.580000 11.845000 -1.400000 13.025000 ;
      RECT -2.580000 13.445000 -1.400000 14.625000 ;
      RECT -2.580000 15.045000 -1.400000 16.225000 ;
      RECT -2.580000 16.645000 -1.400000 17.825000 ;
      RECT -2.580000 18.245000 -1.400000 19.425000 ;
      RECT -2.580000 19.845000 -1.400000 21.025000 ;
      RECT -2.580000 21.445000 -1.400000 22.625000 ;
      RECT -2.580000 23.045000 -1.400000 24.225000 ;
      RECT -2.580000 24.645000 -1.400000 25.825000 ;
      RECT -2.580000 26.245000 -1.400000 27.425000 ;
      RECT -2.580000 27.845000 -1.400000 29.025000 ;
      RECT -2.580000 29.445000 -1.400000 30.625000 ;
      RECT -2.580000 31.045000 -1.400000 32.225000 ;
      RECT -2.580000 32.645000 -1.400000 33.825000 ;
      RECT -2.580000 34.245000 -1.400000 35.425000 ;
      RECT -2.580000 35.845000 -1.400000 37.025000 ;
      RECT -2.580000 37.445000 -1.400000 38.625000 ;
      RECT -2.580000 39.045000 -1.400000 40.225000 ;
      RECT -2.580000 40.645000 -1.400000 41.825000 ;
      RECT -2.580000 42.245000 -1.400000 43.425000 ;
      RECT -2.580000 43.845000 -1.400000 45.025000 ;
      RECT -2.580000 45.445000 -1.400000 46.625000 ;
      RECT -2.580000 47.045000 -1.400000 48.225000 ;
      RECT -2.580000 48.645000 -1.400000 49.825000 ;
      RECT -2.580000 50.245000 -1.400000 51.425000 ;
      RECT -2.580000 51.845000 -1.400000 53.025000 ;
      RECT -2.580000 53.445000 -1.400000 54.625000 ;
      RECT -2.580000 55.045000 -1.400000 56.225000 ;
      RECT -1.035000  2.230000  0.145000  3.410000 ;
      RECT -0.965000 56.660000  0.215000 57.840000 ;
      RECT  0.565000  0.630000  1.745000  1.810000 ;
      RECT  0.635000 58.260000  1.815000 59.440000 ;
      RECT  2.165000 -0.970000  3.345000  0.210000 ;
      RECT  2.235000 59.860000  3.415000 61.040000 ;
      RECT  3.775000 -2.580000  4.955000 -1.400000 ;
      RECT  3.845000 61.400000  5.025000 62.580000 ;
      RECT  5.375000 -2.580000  6.555000 -1.400000 ;
      RECT  5.445000 61.400000  6.625000 62.580000 ;
      RECT  6.975000 -2.580000  8.155000 -1.400000 ;
      RECT  7.045000 61.400000  8.225000 62.580000 ;
      RECT  8.575000 -2.580000  9.755000 -1.400000 ;
      RECT  8.645000 61.400000  9.825000 62.580000 ;
      RECT 10.175000 -2.580000 11.355000 -1.400000 ;
      RECT 10.245000 61.400000 11.425000 62.580000 ;
      RECT 11.775000 -2.580000 12.955000 -1.400000 ;
      RECT 11.845000 61.400000 13.025000 62.580000 ;
      RECT 13.375000 -2.580000 14.555000 -1.400000 ;
      RECT 13.445000 61.400000 14.625000 62.580000 ;
      RECT 14.975000 -2.580000 16.155000 -1.400000 ;
      RECT 15.045000 61.400000 16.225000 62.580000 ;
      RECT 16.575000 -2.580000 17.755000 -1.400000 ;
      RECT 16.645000 61.400000 17.825000 62.580000 ;
      RECT 18.175000 -2.580000 19.355000 -1.400000 ;
      RECT 18.245000 61.400000 19.425000 62.580000 ;
      RECT 19.775000 -2.580000 20.955000 -1.400000 ;
      RECT 19.845000 61.400000 21.025000 62.580000 ;
      RECT 21.375000 -2.580000 22.555000 -1.400000 ;
      RECT 21.445000 61.400000 22.625000 62.580000 ;
      RECT 22.975000 -2.580000 24.155000 -1.400000 ;
      RECT 23.045000 61.400000 24.225000 62.580000 ;
      RECT 24.575000 -2.580000 25.755000 -1.400000 ;
      RECT 24.645000 61.400000 25.825000 62.580000 ;
      RECT 26.175000 -2.580000 27.355000 -1.400000 ;
      RECT 26.245000 61.400000 27.425000 62.580000 ;
      RECT 27.775000 -2.580000 28.955000 -1.400000 ;
      RECT 27.845000 61.400000 29.025000 62.580000 ;
      RECT 29.375000 -2.580000 30.555000 -1.400000 ;
      RECT 29.445000 61.400000 30.625000 62.580000 ;
      RECT 30.975000 -2.580000 32.155000 -1.400000 ;
      RECT 31.045000 61.400000 32.225000 62.580000 ;
      RECT 32.575000 -2.580000 33.755000 -1.400000 ;
      RECT 32.645000 61.400000 33.825000 62.580000 ;
      RECT 34.175000 -2.580000 35.355000 -1.400000 ;
      RECT 34.245000 61.400000 35.425000 62.580000 ;
      RECT 35.775000 -2.580000 36.955000 -1.400000 ;
      RECT 35.845000 61.400000 37.025000 62.580000 ;
      RECT 37.375000 -2.580000 38.555000 -1.400000 ;
      RECT 37.445000 61.400000 38.625000 62.580000 ;
      RECT 38.975000 -2.580000 40.155000 -1.400000 ;
      RECT 39.045000 61.400000 40.225000 62.580000 ;
      RECT 40.575000 -2.580000 41.755000 -1.400000 ;
      RECT 40.645000 61.400000 41.825000 62.580000 ;
      RECT 42.175000 -2.580000 43.355000 -1.400000 ;
      RECT 42.245000 61.400000 43.425000 62.580000 ;
      RECT 43.775000 -2.580000 44.955000 -1.400000 ;
      RECT 43.845000 61.400000 45.025000 62.580000 ;
      RECT 45.375000 -2.580000 46.555000 -1.400000 ;
      RECT 45.445000 61.400000 46.625000 62.580000 ;
      RECT 46.975000 -2.580000 48.155000 -1.400000 ;
      RECT 47.045000 61.400000 48.225000 62.580000 ;
      RECT 48.575000 -2.580000 49.755000 -1.400000 ;
      RECT 48.645000 61.400000 49.825000 62.580000 ;
      RECT 50.175000 -2.580000 51.355000 -1.400000 ;
      RECT 50.245000 61.400000 51.425000 62.580000 ;
      RECT 51.775000 -2.580000 52.955000 -1.400000 ;
      RECT 51.845000 61.400000 53.025000 62.580000 ;
      RECT 53.375000 -2.580000 54.555000 -1.400000 ;
      RECT 53.445000 61.400000 54.625000 62.580000 ;
      RECT 54.975000 -2.580000 56.155000 -1.400000 ;
      RECT 55.045000 61.400000 56.225000 62.580000 ;
      RECT 56.585000 -1.040000 57.765000  0.140000 ;
      RECT 56.655000 59.790000 57.835000 60.970000 ;
      RECT 58.185000  0.560000 59.365000  1.740000 ;
      RECT 58.255000 58.190000 59.435000 59.370000 ;
      RECT 59.785000  2.160000 60.965000  3.340000 ;
      RECT 59.855000 56.590000 61.035000 57.770000 ;
      RECT 61.400000  3.775000 62.580000  4.955000 ;
      RECT 61.400000  5.375000 62.580000  6.555000 ;
      RECT 61.400000  6.975000 62.580000  8.155000 ;
      RECT 61.400000  8.575000 62.580000  9.755000 ;
      RECT 61.400000 10.175000 62.580000 11.355000 ;
      RECT 61.400000 11.775000 62.580000 12.955000 ;
      RECT 61.400000 13.375000 62.580000 14.555000 ;
      RECT 61.400000 14.975000 62.580000 16.155000 ;
      RECT 61.400000 16.575000 62.580000 17.755000 ;
      RECT 61.400000 18.175000 62.580000 19.355000 ;
      RECT 61.400000 19.775000 62.580000 20.955000 ;
      RECT 61.400000 21.375000 62.580000 22.555000 ;
      RECT 61.400000 22.975000 62.580000 24.155000 ;
      RECT 61.400000 24.575000 62.580000 25.755000 ;
      RECT 61.400000 26.175000 62.580000 27.355000 ;
      RECT 61.400000 27.775000 62.580000 28.955000 ;
      RECT 61.400000 29.375000 62.580000 30.555000 ;
      RECT 61.400000 30.975000 62.580000 32.155000 ;
      RECT 61.400000 32.575000 62.580000 33.755000 ;
      RECT 61.400000 34.175000 62.580000 35.355000 ;
      RECT 61.400000 35.775000 62.580000 36.955000 ;
      RECT 61.400000 37.375000 62.580000 38.555000 ;
      RECT 61.400000 38.975000 62.580000 40.155000 ;
      RECT 61.400000 40.575000 62.580000 41.755000 ;
      RECT 61.400000 42.175000 62.580000 43.355000 ;
      RECT 61.400000 43.775000 62.580000 44.955000 ;
      RECT 61.400000 45.375000 62.580000 46.555000 ;
      RECT 61.400000 46.975000 62.580000 48.155000 ;
      RECT 61.400000 48.575000 62.580000 49.755000 ;
      RECT 61.400000 50.175000 62.580000 51.355000 ;
      RECT 61.400000 51.775000 62.580000 52.955000 ;
      RECT 61.400000 53.375000 62.580000 54.555000 ;
      RECT 61.400000 54.975000 62.580000 56.155000 ;
  END
END sky130_fd_pr__padplhp__example_179573804
END LIBRARY
