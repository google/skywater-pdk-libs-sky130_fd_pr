* Copyright 2022 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

******* SkyWater sky130 model library *********
*
* This file is for use by ngspice using the ".lib" statement to select
* a simulation type or corner.  The defined sections are as follows:
*
* Basic corners:
*
* tt  --- Typical N/P device, nominal resistance, nominal capacitance
* ss  --- Slow  N/P device, nominal resistance, nominal capacitance
* sf  --- Slow N/Fast P device, nominal resistance, nominal capacitance
* fs  --- Fast N/Slow P device, nominal resistance, nominal capacitance
* ll  --- Typical N/P device, low resistance, low capacitance
* hl  --- Typical N/P device, high resistance, low capacitance
* lh  --- Typical N/P device, low resistance, high capacitance
* hh  --- Typical N/P device, high resistance, high capacitance
*
* Corners with mismatch analysis:
*
* tt_mm  --- Typical N/P device, nominal resistance, nominal capacitance
* ss_mm  --- Slow  N/P device, nominal resistance, nominal capacitance
* sf_mm  --- Slow N/Fast P device, nominal resistance, nominal capacitance
* fs_mm  --- Fast N/Slow P device, nominal resistance, nominal capacitance
* ll_mm  --- Typical N/P device, low resistance, low capacitance
* hl_mm  --- Typical N/P device, high resistance, low capacitance
* lh_mm  --- Typical N/P device, low resistance, high capacitance
* hh_mm  --- Typical N/P device, high resistance, high capacitance
*
* Monte carlo analysis (process variation):
*
* mc  --- Process Monte Carlo models
*
***********************************************

* Typical corner (tt)
.lib tt
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl tt

* Slow-Fast corner (sf)
.lib sf
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_sf.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl sf

* Fast-Fast corner (ff)
.lib ff
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_ff.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ff

* Slow-Slow corner (ss)
.lib ss
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_ss.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ss

* Fast-Slow corner (fs)
.lib fs
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_fs.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl fs

* Low-Low corner (ll)
.lib ll
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_low.spice
.include parameters_cap_low.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ll

* High-High corner (hh)
.lib hh
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_high.spice
.include parameters_cap_high.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl hh

* High-Low corner (hl)
.lib hl
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_high.spice
.include parameters_cap_low.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl hl

* Low-High corner (lh)
.lib lh
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_low.spice
.include parameters_cap_high.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl lh

* Typical corner with mismatch (tt_mm)
.lib tt_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl tt_mm

* Slow-Fast corner with mismatch (sf_mm)
.lib sf_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_sf.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl sf_mm

* Fast-Fast corner with mismatch (ff_mm)
.lib ff_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_ff.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ff_mm

* Slow-Slow corner with mismatch (ss_mm)
.lib ss_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_ss.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ss_mm

* Fast-Slow corner with mismatch (fs_mm)
.lib fs_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_fs.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl fs_mm

* Low-Low corner with mismatch (ll_mm)
.lib ll_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_low.spice
.include parameters_cap_low.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl ll_mm

* High-High corner with mismatch (hh_mm)
.lib hh_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_high.spice
.include parameters_cap_high.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl hh_mm

* High-Low corner with mismatch (hl_mm)
.lib hl_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_high.spice
.include parameters_cap_low.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl hl_mm

* Low-High corner with mismatch (lh_mm)
.lib lh_mm
.param MC_MM_SWITCH=1
.param MC_PR_SWITCH=0
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_low.spice
.include parameters_cap_high.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl lh_mm

* Monte Carlo process variation
.lib mc
.param MC_MM_SWITCH=0
.param MC_PR_SWITCH=1
.param corner_factor=1
.param process_mc_factor=1
.param mismatch_factor=1

.include parameters_fet_tt.spice
.include parameters_res_nom.spice
.include parameters_cap_nom.spice

* Include the model files
.include models_global.spice
.include models_fet.spice
.include models_bjt.spice
.include models_diodes.spice
.include models_resistors.spice
.include models_capacitors.spice
.endl mc

