# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__pnp_05v5_W3p40L3p40
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pnp_05v5_W3p40L3p40 ;
  ORIGIN -0.130000 -0.130000 ;
  SIZE  6.440000 BY  6.440000 ;
  PIN BASE
    ANTENNADIFFAREA  6.408000 ;
    ANTENNAGATEAREA  26.728899 ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.945000 5.755000 1.305000 ;
        RECT 0.945000 1.305000 1.305000 5.395000 ;
        RECT 0.945000 5.395000 5.755000 5.755000 ;
        RECT 5.395000 1.305000 5.755000 5.395000 ;
    END
  END BASE
  PIN COLLECTOR
    ANTENNADIFFAREA  11.98870 ;
    PORT
      LAYER li1 ;
        RECT 0.130000 0.130000 6.570000 0.625000 ;
        RECT 0.130000 0.625000 0.625000 6.075000 ;
        RECT 0.130000 6.075000 6.570000 6.570000 ;
        RECT 6.075000 0.625000 6.570000 6.075000 ;
    END
  END COLLECTOR
  PIN EMITTER
    ANTENNADIFFAREA  11.559999 ;
    PORT
      LAYER met1 ;
        RECT 1.825000 1.825000 4.875000 4.875000 ;
    END
  END EMITTER
  OBS
    LAYER li1 ;
      RECT 1.615000 1.615000 5.085000 5.085000 ;
    LAYER mcon ;
      RECT 1.980000 1.980000 2.150000 2.150000 ;
      RECT 1.980000 2.480000 2.150000 2.650000 ;
      RECT 1.980000 2.980000 2.150000 3.150000 ;
      RECT 1.980000 3.480000 2.150000 3.650000 ;
      RECT 1.980000 3.980000 2.150000 4.150000 ;
      RECT 1.980000 4.480000 2.150000 4.650000 ;
      RECT 2.480000 1.980000 2.650000 2.150000 ;
      RECT 2.480000 2.480000 2.650000 2.650000 ;
      RECT 2.480000 2.980000 2.650000 3.150000 ;
      RECT 2.480000 3.480000 2.650000 3.650000 ;
      RECT 2.480000 3.980000 2.650000 4.150000 ;
      RECT 2.480000 4.480000 2.650000 4.650000 ;
      RECT 2.980000 1.980000 3.150000 2.150000 ;
      RECT 2.980000 2.480000 3.150000 2.650000 ;
      RECT 2.980000 2.980000 3.150000 3.150000 ;
      RECT 2.980000 3.480000 3.150000 3.650000 ;
      RECT 2.980000 3.980000 3.150000 4.150000 ;
      RECT 2.980000 4.480000 3.150000 4.650000 ;
      RECT 3.480000 1.980000 3.650000 2.150000 ;
      RECT 3.480000 2.480000 3.650000 2.650000 ;
      RECT 3.480000 2.980000 3.650000 3.150000 ;
      RECT 3.480000 3.480000 3.650000 3.650000 ;
      RECT 3.480000 3.980000 3.650000 4.150000 ;
      RECT 3.480000 4.480000 3.650000 4.650000 ;
      RECT 3.980000 1.980000 4.150000 2.150000 ;
      RECT 3.980000 2.480000 4.150000 2.650000 ;
      RECT 3.980000 2.980000 4.150000 3.150000 ;
      RECT 3.980000 3.480000 4.150000 3.650000 ;
      RECT 3.980000 3.980000 4.150000 4.150000 ;
      RECT 3.980000 4.480000 4.150000 4.650000 ;
      RECT 4.480000 1.980000 4.650000 2.150000 ;
      RECT 4.480000 2.480000 4.650000 2.650000 ;
      RECT 4.480000 2.980000 4.650000 3.150000 ;
      RECT 4.480000 3.480000 4.650000 3.650000 ;
      RECT 4.480000 3.980000 4.650000 4.150000 ;
      RECT 4.480000 4.480000 4.650000 4.650000 ;
  END
END sky130_fd_pr__pnp_05v5_W3p40L3p40
END LIBRARY
