* Bipolar transistor I-V characteristic
.param TEMP=27

* Include SkyWater sky130 device models
.include "../../../models/corners/tt/nonfet.spice"
.include "../../../models/sky130_fd_pr__model__pnp.model.spice"

* Base bias
Rb 1 2 680
X1 3 2 5 5 sky130_fd_pr__pnp_05v5_W0p68L0p68 M=1
Rc 3 4 100

* DC source for current measure
Vic 0 4 DC 0V
Vbb 5 1 DC 0V
Vce 5 0 DC 0V

.control
* Sweep Vce from 0 to 1.8V
dc Vce 0 1.8 0.01 Vbb 0 1.2 0.01
let vc1 = V(5) - V(3)
let vb1 = V(5) - V(2)
wrdata sky130_fd_pr__pnp_05v5_W0p68L0p68__iv.data -Vic#branch vb1 vc1

* Sweep Vce from 0 to 3.3V, Vbb from 0 to 2.0V
dc Vce 0 3.3 0.02 Vbb 0.6 0.9 0.01
let beta = Vic#branch / Vbb#branch
let vc2 = V(5) - V(3)
let vb2 = V(5) - V(2)
wrdata sky130_fd_pr__pnp_05v5_W0p68L0p68__beta.data beta vb2 vc2
echo maximum beta
print maximum(beta)
quit
.endc
.end
