# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__res_high_po_0p35__example1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__res_high_po_0p35__example1 ;
  ORIGIN  2.080000  0.000000 ;
  SIZE  4.510000 BY  0.350000 ;
  OBS
    LAYER li1 ;
      RECT -2.080000 0.000000 0.080000 0.350000 ;
      RECT  0.270000 0.000000 2.430000 0.350000 ;
    LAYER mcon ;
      RECT -1.970000 0.090000 -1.800000 0.260000 ;
      RECT -1.610000 0.090000 -1.440000 0.260000 ;
      RECT -1.250000 0.090000 -1.080000 0.260000 ;
      RECT -0.890000 0.090000 -0.720000 0.260000 ;
      RECT -0.530000 0.090000 -0.360000 0.260000 ;
      RECT -0.170000 0.090000  0.000000 0.260000 ;
      RECT  0.350000 0.090000  0.520000 0.260000 ;
      RECT  0.710000 0.090000  0.880000 0.260000 ;
      RECT  1.070000 0.090000  1.240000 0.260000 ;
      RECT  1.430000 0.090000  1.600000 0.260000 ;
      RECT  1.790000 0.090000  1.960000 0.260000 ;
      RECT  2.150000 0.090000  2.320000 0.260000 ;
    LAYER met1 ;
      RECT -2.030000 0.030000 0.060000 0.320000 ;
      RECT  0.290000 0.030000 2.380000 0.320000 ;
  END
END sky130_fd_pr__res_high_po_0p35__example1
END LIBRARY
