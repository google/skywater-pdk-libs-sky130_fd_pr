* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_hvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.255e-06 wmax = 1.265e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.099+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0793014
+ k2 = {-0.20044131+sky130_fd_pr__pfet_01v8_hvt__k2_diff_0}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {83438+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0}
+ ua = {-2.1868798e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_0}
+ ub = {1.7722077e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_0}
+ uc = -1.6417456e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.002956+sky130_fd_pr__pfet_01v8_hvt__u0_diff_0}
+ a0 = {0.65888+sky130_fd_pr__pfet_01v8_hvt__a0_diff_0}
+ keta = {-0.047528+sky130_fd_pr__pfet_01v8_hvt__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.65104277
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_0}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_0}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2637777+sky130_fd_pr__pfet_01v8_hvt__voff_diff_0+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6513386+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.16306432+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0}
+ etab = -0.026662586
+ dsub = 0.35818196
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.72203134+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0}
+ pdiblc1 = 0.38441605
+ pdiblc2 = 0.0078574606
+ pdiblcb = -0.225
+ drout = 0.63135838
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2312485e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.4343701
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.6478246e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.54438+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0}
+ kt2 = -0.053141
+ at = 29266.0
+ ute = -0.279
+ ua1 = 4.3057e-10
+ ub1 = -1.4175e-19
+ uc1 = -5.2391e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.675e-06 wmax = 1.685e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0955+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0888183
+ k2 = {-0.20196049+sky130_fd_pr__pfet_01v8_hvt__k2_diff_1}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {87563+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1}
+ ua = {-2.1838377e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_1}
+ ub = {1.8080364e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_1}
+ uc = -1.1831763e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.003135+sky130_fd_pr__pfet_01v8_hvt__u0_diff_1}
+ a0 = {0.65345+sky130_fd_pr__pfet_01v8_hvt__a0_diff_1}
+ keta = {-0.017748+sky130_fd_pr__pfet_01v8_hvt__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.69867026
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_1}
+ b0 = {2.1073e-024+sky130_fd_pr__pfet_01v8_hvt__b0_diff_1}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24702924+sky130_fd_pr__pfet_01v8_hvt__voff_diff_1+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.15222921+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1}
+ etab = -0.045415713
+ dsub = 0.2958736
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.66659106+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1}
+ pdiblc1 = 0.16607535
+ pdiblc2 = 0.0040091595
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 7.9962646e+8
+ pscbe2 = 7.7649067e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.2550319
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.7051481e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.54438+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1}
+ kt2 = -0.053141
+ at = 29266.0
+ ute = -0.279
+ ua1 = 4.7797e-10
+ ub1 = -1.4175e-19
+ uc1 = -5.2391e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.06+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.51618769
+ k2 = {-0.00083146984+sky130_fd_pr__pfet_01v8_hvt__k2_diff_2}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47380+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2}
+ ua = {-8.5137452e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_2}
+ ub = {6.7844555e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_2}
+ uc = -6.4729555e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0067181+sky130_fd_pr__pfet_01v8_hvt__u0_diff_2}
+ a0 = {0.97582+sky130_fd_pr__pfet_01v8_hvt__a0_diff_2}
+ keta = {-0.013695+sky130_fd_pr__pfet_01v8_hvt__keta_diff_2}
+ a1 = 0.0
+ a2 = 1.0
+ ags = {0.60209+sky130_fd_pr__pfet_01v8_hvt__ags_diff_2}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_2}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16525691+sky130_fd_pr__pfet_01v8_hvt__voff_diff_2+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6996765+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.22+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2}
+ etab = -0.82588402
+ dsub = 0.77677847
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.80609743+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2}
+ pdiblc1 = 0.039
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 7.8630226e+8
+ pscbe2 = 9.1767556e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.6682293
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.0805694e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47906474+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2}
+ kt2 = -0.048559181
+ at = 61761.743
+ ute = -1.0481598
+ ua1 = -4.3040399e-10
+ ub1 = 8.9488555e-19
+ uc1 = 6.6918782e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.09+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43605257
+ k2 = {0.032821892+sky130_fd_pr__pfet_01v8_hvt__k2_diff_3}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53438+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3}
+ ua = {-4.2142258e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_3}
+ ub = {5.0507813e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_3}
+ uc = -6.9850429e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0088976+sky130_fd_pr__pfet_01v8_hvt__u0_diff_3}
+ a0 = {1.1633+sky130_fd_pr__pfet_01v8_hvt__a0_diff_3}
+ keta = {-0.012264+sky130_fd_pr__pfet_01v8_hvt__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.39463+sky130_fd_pr__pfet_01v8_hvt__ags_diff_3}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_3}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17697341+sky130_fd_pr__pfet_01v8_hvt__voff_diff_3+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8787862+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3}
+ etab = -0.00049875119
+ dsub = 0.26129899
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63260008+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.9224047e+8
+ pscbe2 = 9.3515819e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.7757668
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3029923e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46892+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3}
+ kt2 = -0.052362
+ at = 79192.0
+ ute = -0.067643
+ ua1 = 2.8149e-9
+ ub1 = -1.658e-18
+ uc1 = -2.9687e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.085+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43941017
+ k2 = {0.032916976+sky130_fd_pr__pfet_01v8_hvt__k2_diff_4}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53438+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4}
+ ua = {-5.5731408e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_4}
+ ub = {5.6552327e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_4}
+ uc = -7.2710309e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0082748+sky130_fd_pr__pfet_01v8_hvt__u0_diff_4}
+ a0 = {1.1265+sky130_fd_pr__pfet_01v8_hvt__a0_diff_4}
+ keta = {-0.0028979+sky130_fd_pr__pfet_01v8_hvt__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.2984+sky130_fd_pr__pfet_01v8_hvt__ags_diff_4}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_4}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17780505+sky130_fd_pr__pfet_01v8_hvt__voff_diff_4+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2671741+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.041787811+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0020262295
+ pdiblcb = -0.061388807
+ drout = 0.56
+ pscbe1 = 3.7518755e+8
+ pscbe2 = 2.7835156e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.110948
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.9969637e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47523+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4}
+ kt2 = -0.056301
+ at = 90676.0
+ ute = -0.1
+ ua1 = 3.0678e-9
+ ub1 = -2.2467e-18
+ uc1 = -5.8909e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0869+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = {0.03180011+sky130_fd_pr__pfet_01v8_hvt__k2_diff_5}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {160310+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5}
+ ua = {-6.9182204e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_5}
+ ub = {6.2220111e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_5}
+ uc = -7.1776909e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0074657+sky130_fd_pr__pfet_01v8_hvt__u0_diff_5}
+ a0 = {1.2929+sky130_fd_pr__pfet_01v8_hvt__a0_diff_5}
+ keta = {-0.0018702+sky130_fd_pr__pfet_01v8_hvt__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.20339+sky130_fd_pr__pfet_01v8_hvt__ags_diff_5}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_5}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16977492+sky130_fd_pr__pfet_01v8_hvt__voff_diff_5+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5535929+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14095898+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 7.9995125e+8
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.4509773e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5}
+ egidl = 0.88544965
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4407715+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5}
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0779+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0780173
+ k2 = {-0.18691096+sky130_fd_pr__pfet_01v8_hvt__k2_diff_6}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {79622+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6}
+ ua = {-2.368583e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_6}
+ ub = {1.9765955e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_6}
+ uc = 1.6311334e-14
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0024007+sky130_fd_pr__pfet_01v8_hvt__u0_diff_6}
+ a0 = {0.91681+sky130_fd_pr__pfet_01v8_hvt__a0_diff_6}
+ keta = {-0.00052252+sky130_fd_pr__pfet_01v8_hvt__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.80650859
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2174285+sky130_fd_pr__pfet_01v8_hvt__voff_diff_6+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0490306+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.20189086+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6}
+ etab = -0.011570413
+ dsub = 0.30255915
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62222713+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6}
+ pdiblc1 = 0.15311682
+ pdiblc2 = 0.0028344223
+ pdiblcb = -0.3375
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.337696e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.2294593
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.3637136e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.56627+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6}
+ kt2 = -0.096259
+ at = 22259.0
+ ute = -0.005
+ ua1 = 7.4358e-10
+ ub1 = -4.726e-19
+ uc1 = -2.1939e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.042+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.94407842
+ k2 = {-0.14337103+sky130_fd_pr__pfet_01v8_hvt__k2_diff_7}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {104810+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7}
+ ua = {-2.0188743e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_7}
+ ub = {1.650047e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_7}
+ uc = -9.8303269e-12
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0031722+sky130_fd_pr__pfet_01v8_hvt__u0_diff_7}
+ a0 = {0.91559+sky130_fd_pr__pfet_01v8_hvt__a0_diff_7}
+ keta = {-0.050899+sky130_fd_pr__pfet_01v8_hvt__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.5695275
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_7}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_7}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2327165+sky130_fd_pr__pfet_01v8_hvt__voff_diff_7+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.40771457+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7}
+ etab = -6.25e-6
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.68363325+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7}
+ pdiblc1 = 0.39829528
+ pdiblc2 = 0.0099382197
+ pdiblcb = -0.13364569
+ drout = 0.48956724
+ pscbe1 = 8.0e+8
+ pscbe2 = 6.6568323e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.2562888
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.2466963e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53838+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7}
+ kt2 = -0.043005
+ at = 51186.0
+ ute = -0.2477
+ ua1 = 1.9461e-10
+ ub1 = 3.6838e-19
+ uc1 = -3.5153e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0442+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53635572
+ k2 = {0.0035773373+sky130_fd_pr__pfet_01v8_hvt__k2_diff_8}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {99914+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8}
+ ua = {-1.397948e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_8}
+ ub = {1.3291225e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_8}
+ uc = 4.7630651e-14
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0061847+sky130_fd_pr__pfet_01v8_hvt__u0_diff_8}
+ a0 = {0.5931+sky130_fd_pr__pfet_01v8_hvt__a0_diff_8}
+ keta = {-0.033312+sky130_fd_pr__pfet_01v8_hvt__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.5276+sky130_fd_pr__pfet_01v8_hvt__ags_diff_8}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_8}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18912915+sky130_fd_pr__pfet_01v8_hvt__voff_diff_8+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8679711+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8}
+ etab = -6.25e-6
+ dsub = 0.81406049
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63858212+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8}
+ pdiblc1 = 0.40879522
+ pdiblc2 = 0.009193408
+ pdiblcb = -0.21648732
+ drout = 0.48906552
+ pscbe1 = 7.9997105e+8
+ pscbe2 = 9.1548868e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.9566797
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8}
+ bgidl = {1.2603679e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51740568+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8}
+ kt2 = -0.052983574
+ at = 72057.362
+ ute = -0.86411948
+ ua1 = 2.9041801e-10
+ ub1 = -1.7398229e-19
+ uc1 = -1.0365078e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.052+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.516034
+ k2 = {0.0081959434+sky130_fd_pr__pfet_01v8_hvt__k2_diff_9}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55200+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9}
+ ua = {-1.2925874e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_9}
+ ub = {1.0037169e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_9}
+ uc = -2.9729077e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0052584+sky130_fd_pr__pfet_01v8_hvt__u0_diff_9}
+ a0 = {0.71649+sky130_fd_pr__pfet_01v8_hvt__a0_diff_9}
+ keta = {-0.037718+sky130_fd_pr__pfet_01v8_hvt__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.99008978
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_9}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_9}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16535562+sky130_fd_pr__pfet_01v8_hvt__voff_diff_9+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9}
+ etab = -0.000625
+ dsub = 0.26254854
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.027845921+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9}
+ pdiblc1 = 0.011000287
+ pdiblc2 = 4.0135447e-5
+ pdiblcb = -0.019529148
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.32815e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7515738
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.9256988e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53807+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9}
+ kt2 = -0.032665
+ at = 35091.0
+ ute = -0.19855
+ ua1 = 2.5665e-9
+ ub1 = -2.4386e-18
+ uc1 = -1.9533e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0803+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4496415
+ k2 = {0.031927367+sky130_fd_pr__pfet_01v8_hvt__k2_diff_10}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {66641+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10}
+ ua = {-7.3086488e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_10}
+ ub = {6.8083017e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_10}
+ uc = -4.8274863e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0076583+sky130_fd_pr__pfet_01v8_hvt__u0_diff_10}
+ a0 = {1.1973+sky130_fd_pr__pfet_01v8_hvt__a0_diff_10}
+ keta = {-0.014969+sky130_fd_pr__pfet_01v8_hvt__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.57991+sky130_fd_pr__pfet_01v8_hvt__ags_diff_10}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_10}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1661565+sky130_fd_pr__pfet_01v8_hvt__voff_diff_10+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6351533+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.21899552+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10}
+ etab = -0.83278175
+ dsub = 0.73022877
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62281245+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10}
+ pdiblc1 = 0.37098377
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 0.99038333
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2877187e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.8668746
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10}
+ bgidl = {1.2385083e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47253+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10}
+ kt2 = -0.037371
+ at = 102660.0
+ ute = 0.0
+ ua1 = 2.4041e-9
+ ub1 = -1.358e-18
+ uc1 = -9.6365e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0892+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44092059
+ k2 = {0.036899354+sky130_fd_pr__pfet_01v8_hvt__k2_diff_11}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53438+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11}
+ ua = {-3.9144149e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_11}
+ ub = {3.3373675e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_11}
+ uc = -8.5064049e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0083003+sky130_fd_pr__pfet_01v8_hvt__u0_diff_11}
+ a0 = {1.1713+sky130_fd_pr__pfet_01v8_hvt__a0_diff_11}
+ keta = {-0.0087647+sky130_fd_pr__pfet_01v8_hvt__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.3386+sky130_fd_pr__pfet_01v8_hvt__ags_diff_11}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_11}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16593881+sky130_fd_pr__pfet_01v8_hvt__voff_diff_11+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2246948+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33031978+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 2.3783325e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.8248162
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11}
+ bgidl = {1.253884e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.45841675+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11}
+ kt2 = -0.048952895
+ at = 83689.934
+ ute = 0.0
+ ua1 = 2.6153957e-9
+ ub1 = -1.4430041e-18
+ uc1 = 2.893912e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.066+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.51955703
+ k2 = {0.0083255984+sky130_fd_pr__pfet_01v8_hvt__k2_diff_12}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {99197+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12}
+ ua = {-9.2817103e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_12}
+ ub = {6.1068677e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_12}
+ uc = -7.5981588e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0057978+sky130_fd_pr__pfet_01v8_hvt__u0_diff_12}
+ a0 = {1.606+sky130_fd_pr__pfet_01v8_hvt__a0_diff_12}
+ keta = {-0.025019+sky130_fd_pr__pfet_01v8_hvt__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.43619+sky130_fd_pr__pfet_01v8_hvt__ags_diff_12}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_12}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17804625+sky130_fd_pr__pfet_01v8_hvt__voff_diff_12+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1114012+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.6328125+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0026177282
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5686423e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.6922304
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12}
+ bgidl = {1.1982942e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.40079+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12}
+ kt2 = -0.044551
+ at = 179410.0
+ ute = -0.82248
+ ua1 = -3.3779e-10
+ ub1 = 8.7001e-19
+ uc1 = 6.064e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0909+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = {0.018477076+sky130_fd_pr__pfet_01v8_hvt__k2_diff_13}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {160312.5+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13}
+ ua = {-2.7171319e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_13}
+ ub = {1.9996982e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_13}
+ uc = -1.0920239e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0082068126+sky130_fd_pr__pfet_01v8_hvt__u0_diff_13}
+ a0 = {1.6405626+sky130_fd_pr__pfet_01v8_hvt__a0_diff_13}
+ keta = {-0.031235975+sky130_fd_pr__pfet_01v8_hvt__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.44214755+sky130_fd_pr__pfet_01v8_hvt__ags_diff_13}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_13}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17649492+sky130_fd_pr__pfet_01v8_hvt__voff_diff_13+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2740089+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.060146165+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 7.902596e+8
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4593183e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.45554+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13}
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.104+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0855795
+ k2 = {-0.20531331+sky130_fd_pr__pfet_01v8_hvt__k2_diff_14}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {77969+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14}
+ ua = {-2.2584686e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_14}
+ ub = {1.8337483e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_14}
+ uc = -9.8065539e-12
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0029407+sky130_fd_pr__pfet_01v8_hvt__u0_diff_14}
+ a0 = {0.90036+sky130_fd_pr__pfet_01v8_hvt__a0_diff_14}
+ keta = {-0.010637+sky130_fd_pr__pfet_01v8_hvt__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.761054
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_14}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_14}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.23312602+sky130_fd_pr__pfet_01v8_hvt__voff_diff_14+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.21998134+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14}
+ etab = -0.00044348984
+ dsub = 0.2918116
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62863877+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14}
+ pdiblc1 = 0.16025935
+ pdiblc2 = 0.0035027364
+ pdiblcb = -1.1390625
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3001017e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.0394624
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3101263e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53838+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14}
+ kt2 = -0.053141
+ at = 21076.0
+ ute = -0.279
+ ua1 = 4.1797e-10
+ ub1 = -1.4175e-19
+ uc1 = -2.6191e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0669+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.96142823
+ k2 = {-0.14861287+sky130_fd_pr__pfet_01v8_hvt__k2_diff_15}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {85448+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15}
+ ua = {-2.0849956e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_15}
+ ub = {1.6536446e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_15}
+ uc = -8.324554e-12
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0032088+sky130_fd_pr__pfet_01v8_hvt__u0_diff_15}
+ a0 = {0.7581+sky130_fd_pr__pfet_01v8_hvt__a0_diff_15}
+ keta = {-0.073052+sky130_fd_pr__pfet_01v8_hvt__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.66287453
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_15}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_15}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20019295+sky130_fd_pr__pfet_01v8_hvt__voff_diff_15+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8608971+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15}
+ etab = -0.000625
+ dsub = 0.56230341
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.73469042+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15}
+ pdiblc1 = 0.46153647
+ pdiblc2 = 0.0098794151
+ pdiblcb = -0.22461631
+ drout = 0.68441351
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3199817e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.9463947
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.2055002e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51588+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15}
+ kt2 = -0.048792
+ at = 9870.4
+ ute = -0.02
+ ua1 = 8.5338e-10
+ ub1 = -4.6915e-19
+ uc1 = -2.6261e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.04+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.67536437
+ k2 = {-0.053372195+sky130_fd_pr__pfet_01v8_hvt__k2_diff_16}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {82990+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16}
+ ua = {-1.5168868e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_16}
+ ub = {1.2320708e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_16}
+ uc = -1.9527632e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0051814+sky130_fd_pr__pfet_01v8_hvt__u0_diff_16}
+ a0 = {0.7759+sky130_fd_pr__pfet_01v8_hvt__a0_diff_16}
+ keta = {-0.067277+sky130_fd_pr__pfet_01v8_hvt__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {2.2623+sky130_fd_pr__pfet_01v8_hvt__ags_diff_16}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_16}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20169534+sky130_fd_pr__pfet_01v8_hvt__voff_diff_16+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6402517+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16}
+ etab = -0.000625
+ dsub = 0.58604243
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63858582+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16}
+ pdiblc1 = 0.37729626
+ pdiblc2 = 0.0080164025
+ pdiblcb = -0.025
+ drout = 0.43840284
+ pscbe1 = 7.9985266e+8
+ pscbe2 = 9.1408168e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7168788
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16}
+ bgidl = {1.0398522e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.48894097+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16}
+ kt2 = -0.049904433
+ at = 43872.957
+ ute = 0.0
+ ua1 = 1.7802917e-9
+ ub1 = -1.4439577e-18
+ uc1 = -1.173717e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0525+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56908827
+ k2 = {-0.011566694+sky130_fd_pr__pfet_01v8_hvt__k2_diff_17}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {54459+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17}
+ ua = {-1.275487e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_17}
+ ub = {1.0182404e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_17}
+ uc = -3.1964151e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0056349+sky130_fd_pr__pfet_01v8_hvt__u0_diff_17}
+ a0 = {1.1805+sky130_fd_pr__pfet_01v8_hvt__a0_diff_17}
+ keta = {-0.046962+sky130_fd_pr__pfet_01v8_hvt__keta_diff_17}
+ a1 = 0.0
+ a2 = 1.0
+ ags = {1.2529+sky130_fd_pr__pfet_01v8_hvt__ags_diff_17}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_17}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16839389+sky130_fd_pr__pfet_01v8_hvt__voff_diff_17+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6923599+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.076567606+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17}
+ etab = -0.00049978947
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.70967546+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.0010175577
+ pdiblcb = -0.00033376626
+ drout = 0.97122547
+ pscbe1 = 7.9125432e+8
+ pscbe2 = 9.2375409e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.2818518
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17}
+ bgidl = {1.1956507e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.49142+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17}
+ kt2 = -0.047601
+ at = 35000.0
+ ute = -0.02
+ ua1 = 2.1513e-9
+ ub1 = -1.6736e-18
+ uc1 = -7.0232e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0858+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44130134
+ k2 = {0.036889917+sky130_fd_pr__pfet_01v8_hvt__k2_diff_18}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {72710+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18}
+ ua = {-5.3225192e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_18}
+ ub = {5.1388849e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_18}
+ uc = -5.6694956e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0085766+sky130_fd_pr__pfet_01v8_hvt__u0_diff_18}
+ a0 = {1.2006+sky130_fd_pr__pfet_01v8_hvt__a0_diff_18}
+ keta = {-0.013602+sky130_fd_pr__pfet_01v8_hvt__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.54865+sky130_fd_pr__pfet_01v8_hvt__ags_diff_18}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_18}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16518298+sky130_fd_pr__pfet_01v8_hvt__voff_diff_18+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5748567+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.22+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18}
+ etab = -0.30366369
+ dsub = 0.85336401
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60412281+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18}
+ pdiblc1 = 0.38373419
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 0.70261844
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2096545e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.4146004e-5
+ alpha1 = 0.0
+ beta0 = 28.081744
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18}
+ bgidl = {1.3996002e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.48018+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18}
+ kt2 = -0.046569
+ at = 109020.0
+ ute = -1.434
+ ua1 = -3.8899e-10
+ ub1 = 3.2187e-19
+ uc1 = 3.3584e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0872892+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53345147
+ k2 = {0.0027858125+sky130_fd_pr__pfet_01v8_hvt__k2_diff_19}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {35625+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19}
+ ua = {-8.0934302e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_19}
+ ub = {6.7677934e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_19}
+ uc = -5.9955419e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0072052162+sky130_fd_pr__pfet_01v8_hvt__u0_diff_19}
+ a0 = {1.7284184+sky130_fd_pr__pfet_01v8_hvt__a0_diff_19}
+ keta = {-0.063721729+sky130_fd_pr__pfet_01v8_hvt__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.78892655+sky130_fd_pr__pfet_01v8_hvt__ags_diff_19}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_19}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16545197+sky130_fd_pr__pfet_01v8_hvt__voff_diff_19+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1558893+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45648692+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0015421195
+ drout = 0.56
+ pscbe1 = 7.9946973e+8
+ pscbe2 = 9.0633893e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0011084375
+ alpha1 = 0.0
+ beta0 = 34.276539
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19}
+ bgidl = {1.3341834e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.44242368+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19}
+ kt2 = -0.049106631
+ at = 53051.873
+ ute = -0.067525036
+ ua1 = 2.2361689e-9
+ ub1 = -1.259434e-18
+ uc1 = 5.4626174e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0927+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49316523
+ k2 = {0.01697874+sky130_fd_pr__pfet_01v8_hvt__k2_diff_20}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {95427.371+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20}
+ ua = {-3.3723388e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_20}
+ ub = {3.0453411e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_20}
+ uc = -9.1713591e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0086057047+sky130_fd_pr__pfet_01v8_hvt__u0_diff_20}
+ a0 = {1.8+sky130_fd_pr__pfet_01v8_hvt__a0_diff_20}
+ keta = {-0.051588355+sky130_fd_pr__pfet_01v8_hvt__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.60481644+sky130_fd_pr__pfet_01v8_hvt__ags_diff_20}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_20}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1798184+sky130_fd_pr__pfet_01v8_hvt__voff_diff_20+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0684525+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.6328125+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0030509163
+ drout = 0.56
+ pscbe1 = 7.2399674e+8
+ pscbe2 = 9.0530869e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.9685005
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.8443359e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20}
+ bgidl = {2.0270271e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20}
+ egidl = 0.30978258
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.43564+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20}
+ kt2 = -0.044551
+ at = 183070.0
+ ute = -1.192
+ ua1 = -3.3779e-10
+ ub1 = 7.436e-19
+ uc1 = 6.064e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1159+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4341788
+ k2 = {0.038440143+sky130_fd_pr__pfet_01v8_hvt__k2_diff_21}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {160312.5+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21}
+ ua = {-2.1314996e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_21}
+ ub = {4.7411485e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_21}
+ uc = -7.9556859e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.010199256+sky130_fd_pr__pfet_01v8_hvt__u0_diff_21}
+ a0 = {1.665838+sky130_fd_pr__pfet_01v8_hvt__a0_diff_21}
+ keta = {-0.050091678+sky130_fd_pr__pfet_01v8_hvt__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.52002664+sky130_fd_pr__pfet_01v8_hvt__ags_diff_21}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_21}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19418166+sky130_fd_pr__pfet_01v8_hvt__voff_diff_21+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2175692+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.17545984+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00016638736
+ pdiblcb = -0.0030652793
+ drout = 0.56
+ pscbe1 = 7.1874307e+8
+ pscbe2 = 9.6049183e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.7454745e-10
+ alpha1 = 2.7526933e-13
+ beta0 = 3.2147823
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21}
+ bgidl = {1.4504093e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.43169+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21}
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.35073
+ ua1 = 2.2116e-9
+ ub1 = -9.2056e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0954+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0969763
+ k2 = {-0.21116608+sky130_fd_pr__pfet_01v8_hvt__k2_diff_22}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {82498+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22}
+ ua = {-2.2454028e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_22}
+ ub = {1.845539e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_22}
+ uc = -1.0274467e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0031536+sky130_fd_pr__pfet_01v8_hvt__u0_diff_22}
+ a0 = {0.83703+sky130_fd_pr__pfet_01v8_hvt__a0_diff_22}
+ keta = {-0.0081525+sky130_fd_pr__pfet_01v8_hvt__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.79050291
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_22}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_22}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26019244+sky130_fd_pr__pfet_01v8_hvt__voff_diff_22+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.21992699+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22}
+ etab = -0.026458894
+ dsub = 0.29707718
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62670482+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22}
+ pdiblc1 = 0.15132174
+ pdiblc2 = 0.0033763378
+ pdiblcb = -0.253125
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3946251e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.099315
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22}
+ bgidl = {1.0772307e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5204+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22}
+ kt2 = -0.089816
+ at = 44501.0
+ ute = -0.21179
+ ua1 = 1.8804e-10
+ ub1 = 2.6593e-19
+ uc1 = -1.0018e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.096+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.89461406
+ k2 = {-0.13422243+sky130_fd_pr__pfet_01v8_hvt__k2_diff_23}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {102800+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23}
+ ua = {-1.7389301e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_23}
+ ub = {1.3985e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_23}
+ uc = -2.393326e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0046023+sky130_fd_pr__pfet_01v8_hvt__u0_diff_23}
+ a0 = {0.89879+sky130_fd_pr__pfet_01v8_hvt__a0_diff_23}
+ keta = {-0.040629+sky130_fd_pr__pfet_01v8_hvt__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.56974687
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_23}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_23}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.23886342+sky130_fd_pr__pfet_01v8_hvt__voff_diff_23+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.7735611+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23}
+ etab = -0.000625
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.65278044+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23}
+ pdiblc1 = 0.42499332
+ pdiblc2 = 0.0090143058
+ pdiblcb = -0.10470192
+ drout = 0.42008993
+ pscbe1 = 7.9964807e+8
+ pscbe2 = 3.4071835e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.1248308
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23}
+ bgidl = {1.05496e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.48769+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23}
+ kt2 = -0.053086
+ at = 28028.0
+ ute = -0.40375
+ ua1 = 3.7761e-10
+ ub1 = 7.0428e-20
+ uc1 = -9.3567e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.042+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.76036809
+ k2 = {-0.078478762+sky130_fd_pr__pfet_01v8_hvt__k2_diff_24}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {75610+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24}
+ ua = {-1.7682092e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_24}
+ ub = {1.3864375e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_24}
+ uc = -1.3550723e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0045026+sky130_fd_pr__pfet_01v8_hvt__u0_diff_24}
+ a0 = {0.74421+sky130_fd_pr__pfet_01v8_hvt__a0_diff_24}
+ keta = {-0.10038+sky130_fd_pr__pfet_01v8_hvt__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.963+sky130_fd_pr__pfet_01v8_hvt__ags_diff_24}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_24}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20251307+sky130_fd_pr__pfet_01v8_hvt__voff_diff_24+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.490156+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24}
+ etab = -0.000625
+ dsub = 0.7218335
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63775026+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24}
+ pdiblc1 = 0.32127661
+ pdiblc2 = 0.0085305491
+ pdiblcb = -0.025
+ drout = 0.44422126
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.8182288
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24}
+ bgidl = {1.1983673e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47741+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24}
+ kt2 = -0.040182
+ at = 37313.0
+ ute = -0.027
+ ua1 = 1.2301e-9
+ ub1 = -8.8921e-19
+ uc1 = -5.2509e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0644+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4833677
+ k2 = {0.024472177+sky130_fd_pr__pfet_01v8_hvt__k2_diff_25}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {74491+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25}
+ ua = {-1.1805141e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_25}
+ ub = {1.0734439e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_25}
+ uc = -1.0742596e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0067552+sky130_fd_pr__pfet_01v8_hvt__u0_diff_25}
+ a0 = {1.2689+sky130_fd_pr__pfet_01v8_hvt__a0_diff_25}
+ keta = {-0.032245+sky130_fd_pr__pfet_01v8_hvt__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.8312879
+ ags = {1.1009+sky130_fd_pr__pfet_01v8_hvt__ags_diff_25}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_25}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18695718+sky130_fd_pr__pfet_01v8_hvt__voff_diff_25+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4732207+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.054863493+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25}
+ etab = -0.00012499874
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63092942+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25}
+ pdiblc1 = 0.39628238
+ pdiblc2 = 0.0016059821
+ pdiblcb = -0.025
+ drout = 0.70633347
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2926982e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.1501021
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25}
+ bgidl = {1.1645988e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.49132193+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25}
+ kt2 = -0.034228084
+ at = 50649.0
+ ute = -0.11
+ ua1 = 2.5098e-9
+ ub1 = -1.9248e-18
+ uc1 = -1.8195212e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0780308+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4445971
+ k2 = {0.036046509+sky130_fd_pr__pfet_01v8_hvt__k2_diff_26}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {88750.283+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26}
+ ua = {-5.031714e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_26}
+ ub = {4.3050303e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_26}
+ uc = -6.3964987e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0081931334+sky130_fd_pr__pfet_01v8_hvt__u0_diff_26}
+ a0 = {1.8+sky130_fd_pr__pfet_01v8_hvt__a0_diff_26}
+ keta = {-0.041927844+sky130_fd_pr__pfet_01v8_hvt__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.90351153+sky130_fd_pr__pfet_01v8_hvt__ags_diff_26}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_26}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16002206+sky130_fd_pr__pfet_01v8_hvt__voff_diff_26+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.512863+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.21978139+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26}
+ etab = -0.001
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.72200826+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26}
+ pdiblc1 = 0.34455322
+ pdiblc2 = 0.00043
+ pdiblcb = -0.0013402428
+ drout = 0.84940843
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.1042217e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.8119134
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26}
+ bgidl = {1.1265371e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47087793+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26}
+ kt2 = -0.047186161
+ at = 146413.08
+ ute = -1.4106286
+ ua1 = -6.4493406e-10
+ ub1 = 7.6432187e-19
+ uc1 = -2.3969998e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0958+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49484891
+ k2 = {0.016953624+sky130_fd_pr__pfet_01v8_hvt__k2_diff_27}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {56985.594+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27}
+ ua = {-5.0603686e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_27}
+ ub = {4.659009e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_27}
+ uc = -7.278917e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0082826683+sky130_fd_pr__pfet_01v8_hvt__u0_diff_27}
+ a0 = {1.8+sky130_fd_pr__pfet_01v8_hvt__a0_diff_27}
+ keta = {-0.057688775+sky130_fd_pr__pfet_01v8_hvt__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.75329061+sky130_fd_pr__pfet_01v8_hvt__ags_diff_27}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_27}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16625518+sky130_fd_pr__pfet_01v8_hvt__voff_diff_27+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27}
+ etab = -0.0005
+ dsub = 0.35054315
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60908252+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00024386453
+ pdiblcb = -0.0015397845
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6725007e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2919286
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.0527802e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.43067+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27}
+ kt2 = -0.043694
+ at = 90900.0
+ ute = -0.166613
+ ua1 = 1.8352e-9
+ ub1 = -6.365e-19
+ uc1 = -7.2315e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1156+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42968867
+ k2 = {0.039776972+sky130_fd_pr__pfet_01v8_hvt__k2_diff_28}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {125717.43+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28}
+ ua = {-2.0318495e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_28}
+ ub = {5.2559825e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_28}
+ uc = -7.0417557e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.010889942+sky130_fd_pr__pfet_01v8_hvt__u0_diff_28}
+ a0 = {1.8+sky130_fd_pr__pfet_01v8_hvt__a0_diff_28}
+ keta = {-0.055380802+sky130_fd_pr__pfet_01v8_hvt__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.64176685+sky130_fd_pr__pfet_01v8_hvt__ags_diff_28}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_28}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18803206+sky130_fd_pr__pfet_01v8_hvt__voff_diff_28+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2421256+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.6328125+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00047806596
+ pdiblcb = -0.00077107696
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.9505911e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.3164253
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4533856e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.45246+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28}
+ kt2 = -0.040346
+ at = 262510.0
+ ute = -0.29825
+ ua1 = 2.4184e-9
+ ub1 = -9.6782e-19
+ uc1 = 1.3692e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1184+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43657182
+ k2 = {0.038800788+sky130_fd_pr__pfet_01v8_hvt__k2_diff_29}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {200000+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29}
+ ua = {-2.2322697e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_29}
+ ub = {4.8655173e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_29}
+ uc = -7.7670696e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.010379898+sky130_fd_pr__pfet_01v8_hvt__u0_diff_29}
+ a0 = {1.5+sky130_fd_pr__pfet_01v8_hvt__a0_diff_29}
+ keta = {-0.013169082+sky130_fd_pr__pfet_01v8_hvt__keta_diff_29}
+ a1 = 0.0
+ a2 = 1.0
+ ags = {0.3831138+sky130_fd_pr__pfet_01v8_hvt__ags_diff_29}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_29}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18809688+sky130_fd_pr__pfet_01v8_hvt__voff_diff_29+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2739776+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.075489662+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 7.4647513e+8
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29}
+ bgidl = {1.1544446e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.44169+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29}
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0822622
+ k2 = {-0.20530248+sky130_fd_pr__pfet_01v8_hvt__k2_diff_30}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {75665+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30}
+ ua = {-2.2169895e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_30}
+ ub = {1.8138e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_30}
+ uc = -1.5008916e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0033341+sky130_fd_pr__pfet_01v8_hvt__u0_diff_30}
+ a0 = {0.59301+sky130_fd_pr__pfet_01v8_hvt__a0_diff_30}
+ keta = {-0.021696+sky130_fd_pr__pfet_01v8_hvt__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.78383709
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_30}
+ b0 = {2.1073e-024+sky130_fd_pr__pfet_01v8_hvt__b0_diff_30}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.25185386+sky130_fd_pr__pfet_01v8_hvt__voff_diff_30+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.22+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30}
+ etab = -0.035854132
+ dsub = 0.30924623
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62785976+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30}
+ pdiblc1 = 0.17859515
+ pdiblc2 = 0.0038564115
+ pdiblcb = -0.16875
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5148691e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.6340468e-9
+ alpha1 = 0.0
+ beta0 = 13.847471
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30}
+ bgidl = {1.284208e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.52854+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30}
+ kt2 = -0.040578
+ at = 24791.0
+ ute = -0.28
+ ua1 = 4.1289e-10
+ ub1 = -4.1639e-20
+ uc1 = -3.6599e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0638+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.98410246
+ k2 = {-0.15921092+sky130_fd_pr__pfet_01v8_hvt__k2_diff_31}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {75326+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31}
+ ua = {-2.1424017e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_31}
+ ub = {1.6755e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_31}
+ uc = -1.093974e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0032452+sky130_fd_pr__pfet_01v8_hvt__u0_diff_31}
+ a0 = {0.60495+sky130_fd_pr__pfet_01v8_hvt__a0_diff_31}
+ keta = {-0.088216+sky130_fd_pr__pfet_01v8_hvt__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.7245882
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_31}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_31}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2086929+sky130_fd_pr__pfet_01v8_hvt__voff_diff_31+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6948856+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31}
+ etab = -0.00062500003
+ dsub = 0.56499453
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.70320506+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31}
+ pdiblc1 = 0.40758103
+ pdiblc2 = 0.0091365927
+ pdiblcb = -0.17539027
+ drout = 0.58508493
+ pscbe1 = 7.9989774e+8
+ pscbe2 = 9.2821999e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.4511866e-8
+ alpha1 = 0.0
+ beta0 = 16.184805
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31}
+ bgidl = {1.397257e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31}
+ cgidl = {49.03999+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51769+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31}
+ kt2 = -0.053086
+ at = 33028.0
+ ute = -0.16694
+ ua1 = 3.7761e-10
+ ub1 = 7.0428e-20
+ uc1 = -9.3567e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.056+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.7471885
+ k2 = {-0.07475736+sky130_fd_pr__pfet_01v8_hvt__k2_diff_32}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {81648+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32}
+ ua = {-1.8602371e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_32}
+ ub = {1.5376e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_32}
+ uc = 2.0393181e-14
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0046393+sky130_fd_pr__pfet_01v8_hvt__u0_diff_32}
+ a0 = {0.78195+sky130_fd_pr__pfet_01v8_hvt__a0_diff_32}
+ keta = {-0.087499+sky130_fd_pr__pfet_01v8_hvt__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {2.3062+sky130_fd_pr__pfet_01v8_hvt__ags_diff_32}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_32}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19332381+sky130_fd_pr__pfet_01v8_hvt__voff_diff_32+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.7961467+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32}
+ etab = -0.000625
+ dsub = 0.68351845
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.72217021+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32}
+ pdiblc1 = 0.37481283
+ pdiblc2 = 0.00847069
+ pdiblcb = -0.025
+ drout = 0.56215143
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.5780878e-8
+ alpha1 = 0.0
+ beta0 = 16.648985
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32}
+ bgidl = {1.2422931e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.49688692+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32}
+ kt2 = -0.038371627
+ at = 45286.948
+ ute = -0.05
+ ua1 = 1.2030437e-9
+ ub1 = -7.4291142e-19
+ uc1 = -7.4139789e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.062+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47940167
+ k2 = {0.025228682+sky130_fd_pr__pfet_01v8_hvt__k2_diff_33}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {76181+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33}
+ ua = {-1.1418974e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_33}
+ ub = {1.0181e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_33}
+ uc = -1.4888633e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0067018+sky130_fd_pr__pfet_01v8_hvt__u0_diff_33}
+ a0 = {1.0839+sky130_fd_pr__pfet_01v8_hvt__a0_diff_33}
+ keta = {-0.030761+sky130_fd_pr__pfet_01v8_hvt__keta_diff_33}
+ a1 = 0.0
+ a2 = 1.0
+ ags = {0.93515+sky130_fd_pr__pfet_01v8_hvt__ags_diff_33}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_33}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17869917+sky130_fd_pr__pfet_01v8_hvt__voff_diff_33+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5089649+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.014184772+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33}
+ etab = -0.001
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.88914551+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33}
+ pdiblc1 = 0.055790472
+ pdiblc2 = 0.00077664689
+ pdiblcb = -0.025
+ drout = 0.9532331
+ pscbe1 = 7.5896555e+8
+ pscbe2 = 9.1354199e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0699549
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33}
+ bgidl = {1.1691122e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4903768+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33}
+ kt2 = -0.032665077
+ at = 40000.0
+ ute = -0.11
+ ua1 = 2.5665e-9
+ ub1 = -2.0842e-18
+ uc1 = -1.9532902e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.48072746
+ k2 = {0.012321803+sky130_fd_pr__pfet_01v8_hvt__k2_diff_34}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {40253+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34}
+ ua = {-1.2162698e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_34}
+ ub = {9.0906101e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_34}
+ uc = -5.3977149e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0062058+sky130_fd_pr__pfet_01v8_hvt__u0_diff_34}
+ a0 = {1.1296+sky130_fd_pr__pfet_01v8_hvt__a0_diff_34}
+ keta = {-0.013884019+sky130_fd_pr__pfet_01v8_hvt__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.80322+sky130_fd_pr__pfet_01v8_hvt__ags_diff_34}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_34}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.15239965+sky130_fd_pr__pfet_01v8_hvt__voff_diff_34+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3341073+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.22+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34}
+ etab = -0.84636554
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.4019278+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34}
+ pdiblc1 = 0.38864941
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.8447626
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.0954252e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.6893915e-11
+ alpha1 = -1.0e-10
+ beta0 = 6.2607413
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.0937505e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46303+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34}
+ kt2 = -0.051385
+ at = 39763.0
+ ute = -1.0096
+ ua1 = -6.0791e-10
+ ub1 = 1.1586e-18
+ uc1 = 1.0712e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0822+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = {0.036341026+sky130_fd_pr__pfet_01v8_hvt__k2_diff_35}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80156+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35}
+ ua = {-6.0301916e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_35}
+ ub = {4.3041395e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_35}
+ uc = -1.0566299e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0074557+sky130_fd_pr__pfet_01v8_hvt__u0_diff_35}
+ a0 = {1.464+sky130_fd_pr__pfet_01v8_hvt__a0_diff_35}
+ keta = {0.023361259+sky130_fd_pr__pfet_01v8_hvt__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.97
+ ags = {0.11329+sky130_fd_pr__pfet_01v8_hvt__ags_diff_35}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_35}
+ b1 = {2.1073e-024+sky130_fd_pr__pfet_01v8_hvt__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17508072+sky130_fd_pr__pfet_01v8_hvt__voff_diff_35+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6473612+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35}
+ cit = 3.2465718e-7
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.015+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.9002574e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.43825+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35}
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0867333+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47183665
+ k2 = {0.018908449+sky130_fd_pr__pfet_01v8_hvt__k2_diff_36}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {50706.805+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36}
+ ua = {-1.0534351e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_36}
+ ub = {7.3416654e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_36}
+ uc = -6.9057193e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0064899791+sky130_fd_pr__pfet_01v8_hvt__u0_diff_36}
+ a0 = {1.2296686+sky130_fd_pr__pfet_01v8_hvt__a0_diff_36}
+ keta = {-0.0010722962+sky130_fd_pr__pfet_01v8_hvt__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.27979705+sky130_fd_pr__pfet_01v8_hvt__ags_diff_36}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_36}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.15888314+sky130_fd_pr__pfet_01v8_hvt__voff_diff_36+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6747976+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36}
+ etab = -0.0005
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63484294+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3781415e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6177381
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.9586586e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53604+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36}
+ kt2 = -0.05223
+ at = 10000.0
+ ute = -1.0659
+ ua1 = 4.5568e-10
+ ub1 = -2.7217e-19
+ uc1 = 5.2142e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.1027+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42180358
+ k2 = {0.034434574+sky130_fd_pr__pfet_01v8_hvt__k2_diff_37}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {54812.074+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37}
+ ua = {-4.5085882e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_37}
+ ub = {3.2682605e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_37}
+ uc = -1.0711711e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0085984431+sky130_fd_pr__pfet_01v8_hvt__u0_diff_37}
+ a0 = {1.2594348+sky130_fd_pr__pfet_01v8_hvt__a0_diff_37}
+ keta = {0.013644534+sky130_fd_pr__pfet_01v8_hvt__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.19308737+sky130_fd_pr__pfet_01v8_hvt__ags_diff_37}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_37}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17662052+sky130_fd_pr__pfet_01v8_hvt__voff_diff_37+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.701106+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.34304825+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00057854717
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5516009e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4740645e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.41825+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37}
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.12298
+ ua1 = 2.0902e-9
+ ub1 = -1.1289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.081+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43148777
+ k2 = {0.033864949+sky130_fd_pr__pfet_01v8_hvt__k2_diff_38}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80156+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38}
+ ua = {-5.3845529e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_38}
+ ub = {3.5204569e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_38}
+ uc = -1.0990767e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0077695+sky130_fd_pr__pfet_01v8_hvt__u0_diff_38}
+ a0 = {1.3962+sky130_fd_pr__pfet_01v8_hvt__a0_diff_38}
+ keta = {0.024383441+sky130_fd_pr__pfet_01v8_hvt__keta_diff_38}
+ a1 = 0.0
+ a2 = 0.97
+ ags = {0.12567+sky130_fd_pr__pfet_01v8_hvt__ags_diff_38}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_38}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_38}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17742247+sky130_fd_pr__pfet_01v8_hvt__voff_diff_38+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4425849+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.017402344+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030866885
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 6.6004928e+8
+ pscbe2 = 9.7083071e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.5013384e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50604+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38}
+ kt2 = -0.05223
+ at = 10000.0
+ ute = -1.0359
+ ua1 = 4.8568e-10
+ ub1 = -2.7217e-19
+ uc1 = 5.2142e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.114+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.97201195
+ k2 = {-0.19535474+sky130_fd_pr__pfet_01v8_hvt__k2_diff_39}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109040+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39}
+ ua = {-2.1578101e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_39}
+ ub = {1.8047023e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_39}
+ uc = -1.9161134e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0031373+sky130_fd_pr__pfet_01v8_hvt__u0_diff_39}
+ a0 = {1.0049776+sky130_fd_pr__pfet_01v8_hvt__a0_diff_39}
+ keta = {-0.017237009+sky130_fd_pr__pfet_01v8_hvt__keta_diff_39}
+ a1 = 0.0
+ a2 = 0.63412408
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_39}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_39}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_39}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19529487+sky130_fd_pr__pfet_01v8_hvt__voff_diff_39+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39}
+ etab = -0.000625
+ dsub = 0.48688771
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62457134+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39}
+ pdiblc1 = 0.16324552
+ pdiblc2 = 0.0037058195
+ pdiblcb = -0.50625
+ drout = 1.0
+ pscbe1 = 7.9999957e+8
+ pscbe2 = 9.4716968e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3819491
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.1396435e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.52214+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39}
+ kt2 = -0.048777
+ at = 37150.0
+ ute = -0.1632
+ ua1 = 8.4379e-10
+ ub1 = -6.2949e-19
+ uc1 = -8.2789e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0764+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.85164386
+ k2 = {-0.12683+sky130_fd_pr__pfet_01v8_hvt__k2_diff_40}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {132400+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40}
+ ua = {-2.164253e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_40}
+ ub = {1.8572189e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_40}
+ uc = 2.58041e-13
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0030964+sky130_fd_pr__pfet_01v8_hvt__u0_diff_40}
+ a0 = {1.166315+sky130_fd_pr__pfet_01v8_hvt__a0_diff_40}
+ keta = {-0.028218739+sky130_fd_pr__pfet_01v8_hvt__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.45249595
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_40}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_40}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18676697+sky130_fd_pr__pfet_01v8_hvt__voff_diff_40+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8760044+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40}
+ etab = -6.25e-6
+ dsub = 0.66213569
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.82665932+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40}
+ pdiblc1 = 0.18776805
+ pdiblc2 = 0.0066944085
+ pdiblcb = -0.225
+ drout = 0.9981043
+ pscbe1 = 7.9996855e+8
+ pscbe2 = 9.3174823e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0852145
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.9262738e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.54112+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40}
+ kt2 = -0.042333
+ at = 105041.0
+ ute = -0.42503
+ ua1 = 2.9333e-10
+ ub1 = 5.4574e-20
+ uc1 = -5.8335e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.119+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50013358
+ k2 = {0.017366908+sky130_fd_pr__pfet_01v8_hvt__k2_diff_41}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {92665+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41}
+ ua = {-1.5575025e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_41}
+ ub = {1.2428657e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_41}
+ uc = -1.7540731e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0051179+sky130_fd_pr__pfet_01v8_hvt__u0_diff_41}
+ a0 = {0.84229689+sky130_fd_pr__pfet_01v8_hvt__a0_diff_41}
+ keta = {-0.02917043+sky130_fd_pr__pfet_01v8_hvt__keta_diff_41}
+ a1 = 0.0
+ a2 = 0.97
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_41}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_41}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_41}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1619475+sky130_fd_pr__pfet_01v8_hvt__voff_diff_41+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8525471+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41}
+ etab = -6.25e-6
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.038924225+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41}
+ pdiblc1 = 0.013035351
+ pdiblc2 = 2.6875e-5
+ pdiblcb = -0.10009403
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.1480723e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.166112
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.9962149e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50388+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41}
+ kt2 = -0.059544
+ at = 80000.0
+ ute = -0.1686
+ ua1 = 1.3219e-9
+ ub1 = -7.9801e-19
+ uc1 = -6.7349e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.066397+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50802186
+ k2 = {0.00893704+sky130_fd_pr__pfet_01v8_hvt__k2_diff_42}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {51812.515+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42}
+ ua = {-1.4244083e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_42}
+ ub = {1.0216384e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_42}
+ uc = -4.3585047e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0048447295+sky130_fd_pr__pfet_01v8_hvt__u0_diff_42}
+ a0 = {1.2572312+sky130_fd_pr__pfet_01v8_hvt__a0_diff_42}
+ keta = {-0.0010368697+sky130_fd_pr__pfet_01v8_hvt__keta_diff_42}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.56427018+sky130_fd_pr__pfet_01v8_hvt__ags_diff_42}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_42}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_42}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.14904922+sky130_fd_pr__pfet_01v8_hvt__voff_diff_42+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4353498+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42}
+ etab = -0.0012469733
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62805205+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42}
+ pdiblc1 = 0.38433914
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.73636547
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.1701202e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.4713014
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.2341059e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47906474+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42}
+ kt2 = -0.048559181
+ at = 51761.743
+ ute = -1.0481598
+ ua1 = -4.3040399e-10
+ ub1 = 8.5488555e-19
+ uc1 = 6.6918782e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0982+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.5072526
+ k2 = {0.00063343074+sky130_fd_pr__pfet_01v8_hvt__k2_diff_43}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {33805+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43}
+ ua = {-7.7290065e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_43}
+ ub = {6.2039968e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_43}
+ uc = -8.117396e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0078733+sky130_fd_pr__pfet_01v8_hvt__u0_diff_43}
+ a0 = {1.1454+sky130_fd_pr__pfet_01v8_hvt__a0_diff_43}
+ keta = {-0.0091786+sky130_fd_pr__pfet_01v8_hvt__keta_diff_43}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.40776+sky130_fd_pr__pfet_01v8_hvt__ags_diff_43}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_43}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_43}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16843277+sky130_fd_pr__pfet_01v8_hvt__voff_diff_43+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8440334+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43}
+ etab = -0.0005
+ dsub = 0.26000001
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.77228851+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00044132367
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4663397e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.5678953
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.2771072e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.45287+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43}
+ kt2 = -0.053935
+ at = 40042.0
+ ute = -0.27335
+ ua1 = 1.3027e-9
+ ub1 = -3.62e-19
+ uc1 = 3.5526e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0928+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44665324
+ k2 = {0.023922352+sky130_fd_pr__pfet_01v8_hvt__k2_diff_44}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {58700.889+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44}
+ ua = {-3.9411538e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_44}
+ ub = {3.4511372e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_44}
+ uc = -1.0733757e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.008771213+sky130_fd_pr__pfet_01v8_hvt__u0_diff_44}
+ a0 = {1.2723362+sky130_fd_pr__pfet_01v8_hvt__a0_diff_44}
+ keta = {0.0067226692+sky130_fd_pr__pfet_01v8_hvt__keta_diff_44}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.18304086+sky130_fd_pr__pfet_01v8_hvt__ags_diff_44}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_44}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_44}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16990138+sky130_fd_pr__pfet_01v8_hvt__voff_diff_44+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.68962544+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.0916125e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.7974328e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.44425+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44}
+ kt2 = -0.058546
+ at = 100990.0
+ ute = -0.18298
+ ua1 = 2.0902e-9
+ ub1 = -1.1289e-18
+ uc1 = -4.1814e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0906866+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.45351162
+ k2 = {0.024555927+sky130_fd_pr__pfet_01v8_hvt__k2_diff_45}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {61064.004+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45}
+ ua = {-4.9723649e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_45}
+ ub = {4.0294943e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_45}
+ uc = -1.0717282e-10
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.008070795+sky130_fd_pr__pfet_01v8_hvt__u0_diff_45}
+ a0 = {1.2209207+sky130_fd_pr__pfet_01v8_hvt__a0_diff_45}
+ keta = {0.0071303363+sky130_fd_pr__pfet_01v8_hvt__keta_diff_45}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.11410703+sky130_fd_pr__pfet_01v8_hvt__ags_diff_45}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_45}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_45}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18613842+sky130_fd_pr__pfet_01v8_hvt__voff_diff_45+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3987334+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14095898+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00033122306
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.1855131e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.3672742e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.42906474+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45}
+ kt2 = -0.048559181
+ at = 61761.743
+ ute = -1.0481598
+ ua1 = -4.3040399e-10
+ ub1 = 8.9488555e-19
+ uc1 = 6.6918782e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0597+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0502231
+ k2 = {-0.18874213+sky130_fd_pr__pfet_01v8_hvt__k2_diff_46}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {85231+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46}
+ ua = {-2.3441206e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_46}
+ ub = {2.0170582e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_46}
+ uc = 1.9113717e-14
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.002497+sky130_fd_pr__pfet_01v8_hvt__u0_diff_46}
+ a0 = {1.0132+sky130_fd_pr__pfet_01v8_hvt__a0_diff_46}
+ keta = {0.04103419+sky130_fd_pr__pfet_01v8_hvt__keta_diff_46}
+ a1 = 0.0
+ a2 = 0.95671944
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_46}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_46}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_46}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.25024889+sky130_fd_pr__pfet_01v8_hvt__voff_diff_46+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6818969+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.18519279+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46}
+ etab = -0.018159526
+ dsub = 0.28488048
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62190714+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46}
+ pdiblc1 = 0.17199343
+ pdiblc2 = 0.0021176917
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 7.8075686e+8
+ pscbe2 = 9.1842717e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.9923957
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.0698583e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.57223+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46}
+ kt2 = -0.093165
+ at = 55755.0
+ ute = -0.1632
+ ua1 = 7.4358e-10
+ ub1 = -6.474e-19
+ uc1 = -4.1394e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.176e-008+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.087+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4349469
+ k2 = {0.033033416+sky130_fd_pr__pfet_01v8_hvt__k2_diff_47}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109430+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47}
+ ua = {-7.9553952e-010+sky130_fd_pr__pfet_01v8_hvt__ua_diff_47}
+ ub = {6.7360576e-019+sky130_fd_pr__pfet_01v8_hvt__ub_diff_47}
+ uc = -4.8332508e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0076558+sky130_fd_pr__pfet_01v8_hvt__u0_diff_47}
+ a0 = {1.1143+sky130_fd_pr__pfet_01v8_hvt__a0_diff_47}
+ keta = {-0.043531+sky130_fd_pr__pfet_01v8_hvt__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.49215603
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_47}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_47}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.16857953+sky130_fd_pr__pfet_01v8_hvt__voff_diff_47+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4777762+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0081705343+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47}
+ etab = -0.00099999893
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.4325064+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47}
+ pdiblc1 = 0.069872306
+ pdiblc2 = 0.00080363033
+ pdiblcb = -0.225
+ drout = 0.51197505
+ pscbe1 = 1.3828473e+8
+ pscbe2 = 7.8174856e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.4421206
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.133969e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.48388+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47}
+ kt2 = -0.059544
+ at = 80000.0
+ ute = -0.2386
+ ua1 = 1.6656e-9
+ ub1 = -8.6644e-19
+ uc1 = -6.7349e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.089+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.0716985
+ k2 = {-0.20271345+sky130_fd_pr__pfet_01v8_hvt__k2_diff_48}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {78922+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48}
+ ua = {-2.2873261e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_48}
+ ub = {1.8906205e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_48}
+ uc = -1.3332403e-11
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.002687+sky130_fd_pr__pfet_01v8_hvt__u0_diff_48}
+ a0 = {0.87713+sky130_fd_pr__pfet_01v8_hvt__a0_diff_48}
+ keta = {-0.012556+sky130_fd_pr__pfet_01v8_hvt__keta_diff_48}
+ a1 = 0.0
+ a2 = 0.74869385
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_48}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_48}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_48}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2025646+sky130_fd_pr__pfet_01v8_hvt__voff_diff_48+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4131397+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48}
+ etab = -0.0008517151
+ dsub = 0.4339823
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62077198+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48}
+ pdiblc1 = 0.35507256
+ pdiblc2 = 0.0012371251
+ pdiblcb = -1.1390625
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 5.1545636e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.353946
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.035337e-009+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.58669+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48}
+ kt2 = -0.050786
+ at = 18280.0
+ ute = -0.48325
+ ua1 = 3.4998e-10
+ ub1 = -1.1387e-19
+ uc1 = -2.9301e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {9.364e-009+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -6.0e-8
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.118+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.1107151
+ k2 = {-0.21107143+sky130_fd_pr__pfet_01v8_hvt__k2_diff_49}
+ k3 = -13.778
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {87856+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49}
+ ua = {-2.3304507e-009+sky130_fd_pr__pfet_01v8_hvt__ua_diff_49}
+ ub = {1.9668119e-018+sky130_fd_pr__pfet_01v8_hvt__ub_diff_49}
+ uc = 8.5835281e-14
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49}
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
+ u0 = {0.0026289+sky130_fd_pr__pfet_01v8_hvt__u0_diff_49}
+ a0 = {1.1333+sky130_fd_pr__pfet_01v8_hvt__a0_diff_49}
+ keta = {0.00077411+sky130_fd_pr__pfet_01v8_hvt__keta_diff_49}
+ a1 = 0.0
+ a2 = 0.64520655
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_49}
+ b0 = {0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_49}
+ b1 = {0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_49}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20169156+sky130_fd_pr__pfet_01v8_hvt__voff_diff_49+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8349351+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.21948109+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49}
+ etab = -0.027368442
+ dsub = 0.30975235
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62207689+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49}
+ pdiblc1 = 0.1677304
+ pdiblc2 = 0.0038590567
+ pdiblcb = -0.3796875
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 7.3782091e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3514574
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.2929704e-010+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49}
+ cgidl = {300+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53627+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49}
+ kt2 = -0.096259
+ at = 41259.0
+ ute = -0.05
+ ua1 = 7.4358e-10
+ ub1 = -4.726e-19
+ uc1 = -2.1939e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2556
+ jss = 2.17e-5
+ jsws = 8.200000000000001e-10
+ xtis = 2.0
+ bvs = 12.8
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0019551
+ tpbsw = 0.00014242
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.0
+ tcjswg = 2.0e-12
+ cgdo = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgso = {6e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdl = {7.6e-012*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.2435e-011*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbsws = 0.7418
+ cjswgs = {2.4701e-010*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
+ pbswgs = 1.3925
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = .0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = .25e-6
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = .25e-6
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos
* Model Flag Parameters
+ lmin = 1.79e-07 lmax = 1.81e-07 wmin = 6.39e-07 wmax = 6.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07095600111241+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.07169844263695
+ k2 = {-0.211129143952937+sky130_fd_pr__pfet_01v8_hvt__k2_diff_50}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.433982266549591
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.294825592439786+sky130_fd_pr__pfet_01v8_hvt__voff_diff_50+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.2192092567159+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.490000000445447+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50}
+ etab = -0.000851725200424369
+ u0 = {0.00265505728828512+sky130_fd_pr__pfet_01v8_hvt__u0_diff_50}
+ ua = {-2.37404714270393e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_50}
+ ub = {2.05009051203083e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_50}
+ uc = -1.33324015760675e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {84343.5987161124+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50}
+ a0 = {0.877130207986808+sky130_fd_pr__pfet_01v8_hvt__a0_diff_50}
+ ags = {1.25000000856918+sky130_fd_pr__pfet_01v8_hvt__ags_diff_50}
+ a1 = 0.0
+ a2 = 0.748693858171036
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_50}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_50}
+ keta = {-0.0125559961514956+sky130_fd_pr__pfet_01v8_hvt__keta_diff_50}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.620771983425462+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50}
+ pdiblc1 = 0.355072622104209
+ pdiblc2 = 0.00123712400757925
+ pdiblcb = -1.13906250407908
+ drout = 1.00000002589623
+ pscbe1 = 800000000.056997
+ pscbe2 = 5.1545629766385e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35394585616203
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {1.03533670551374e-09+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50}
+ bgidl = {1000000043.63208+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.586690043055798+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50}
+ kt2 = -0.0507860334352673
+ at = 18280.0055530857
+ ute = -0.483250041537429
+ ua1 = 3.49980190249352e-10
+ ub1 = -1.13870110915159e-19
+ uc1 = -2.93009994723167e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 1.999e-06 wmax = 2.001e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07847201664917+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.08557951889565
+ k2 = {-0.216553287031283+sky130_fd_pr__pfet_01v8_hvt__k2_diff_51}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.291811607936174
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.274450017810204+sky130_fd_pr__pfet_01v8_hvt__voff_diff_51+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.18742003558682+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.219981332437539+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51}
+ etab = -0.000443489865924838
+ u0 = {0.00332799993611169+sky130_fd_pr__pfet_01v8_hvt__u0_diff_51}
+ ua = {-2.2206406139198e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_51}
+ ub = {1.90440730167961e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_51}
+ uc = -9.80655408020155e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {67715.0255112324+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51}
+ a0 = {0.900359976212471+sky130_fd_pr__pfet_01v8_hvt__a0_diff_51}
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_51}
+ a1 = 0.0
+ a2 = 0.761053992788159
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_51}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_51}
+ keta = {-0.0106370129267269+sky130_fd_pr__pfet_01v8_hvt__keta_diff_51}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.628638745580517+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51}
+ pdiblc1 = 0.160259391056057
+ pdiblc2 = 0.0035027346670166
+ pdiblcb = -1.13906214402687
+ drout = 0.999999942221289
+ pscbe1 = 800000000.0
+ pscbe2 = 9.30010169804745e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.03946235626706
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {1.31012667814403e-10+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51}
+ bgidl = {1000000000.0+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.538380001312198+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51}
+ kt2 = -0.0531410025950031
+ at = 21075.9960193155
+ ute = -0.2789999847785
+ ua1 = 4.17969968549234e-10
+ ub1 = -1.41749973441109e-19
+ uc1 = -2.61909999842536e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 1.119e-06 wmax = 1.121e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07810236233414+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.07801730927071
+ k2 = {-0.21237395755418+sky130_fd_pr__pfet_01v8_hvt__k2_diff_52}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.302559137958808
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.298266481655818+sky130_fd_pr__pfet_01v8_hvt__voff_diff_52+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.18013117522574+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.201890675816754+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52}
+ etab = -0.0115703919135681
+ u0 = {0.00360890031315458+sky130_fd_pr__pfet_01v8_hvt__u0_diff_52}
+ ua = {-2.02168292270409e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_52}
+ ub = {1.73435492221335e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_52}
+ uc = 1.63174963510485e-14
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {78561.9811960684+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52}
+ a0 = {0.91681021358675+sky130_fd_pr__pfet_01v8_hvt__a0_diff_52}
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_52}
+ a1 = 0.0
+ a2 = 0.8065085362853
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_52}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_52}
+ keta = {-0.000522512448261736+sky130_fd_pr__pfet_01v8_hvt__keta_diff_52}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.622227158030407+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52}
+ pdiblc1 = 0.153116553170111
+ pdiblc2 = 0.00283442620341279
+ pdiblcb = -0.33749917040476
+ drout = 1.00000079909858
+ pscbe1 = 800000000.0
+ pscbe2 = 8.3376919564349e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.22945978680628
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {5.36378173239407e-10+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52}
+ bgidl = {1000000000.0+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.5662699807296+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52}
+ kt2 = -0.0962589671051477
+ at = 22258.9879460876
+ ute = -0.00500007502147426
+ ua1 = 7.43579433877174e-10
+ ub1 = -4.72599350433354e-19
+ uc1 = -2.19389545270368e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 1.649e-06 wmax = 1.651e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.08357901503254+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.08881830915389
+ k2 = {-0.218252474805795+sky130_fd_pr__pfet_01v8_hvt__k2_diff_53}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.295873540877598
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.279273238442158+sky130_fd_pr__pfet_01v8_hvt__voff_diff_53+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.50857000762125+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.152229183476801+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53}
+ etab = -0.0454157070816712
+ u0 = {0.00420239993275247+sky130_fd_pr__pfet_01v8_hvt__u0_diff_53}
+ ua = {-1.83797766294352e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_53}
+ ub = {1.5790164508923e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_53}
+ uc = -1.18317630978375e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {80136.1961431871+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53}
+ a0 = {0.653449991929456+sky130_fd_pr__pfet_01v8_hvt__a0_diff_53}
+ ags = {1.25+sky130_fd_pr__pfet_01v8_hvt__ags_diff_53}
+ a1 = 0.0
+ a2 = 0.698670227892085
+ b0 = {2.10730023619567e-24+sky130_fd_pr__pfet_01v8_hvt__b0_diff_53}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_53}
+ keta = {-0.017747994973756+sky130_fd_pr__pfet_01v8_hvt__keta_diff_53}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.666591065931766+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53}
+ pdiblc1 = 0.166075379298761
+ pdiblc2 = 0.00400915914297712
+ pdiblcb = -0.0750000013226959
+ drout = 0.999999942221289
+ pscbe1 = 799626457.465883
+ pscbe2 = 7.76490646951502e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.25503194584925
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {6.70514827923578e-10+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53}
+ bgidl = {1000000000.0+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.544379998162922+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53}
+ kt2 = -0.0531410025950031
+ at = 29266.0042263279
+ ute = -0.2789999847785
+ ua1 = 4.77969989544405e-10
+ ub1 = -1.41749973441109e-19
+ uc1 = -5.23910049842536e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos
* Model Flag Parameters
+ lmin = 1.79e-07 lmax = 1.81e-07 wmin = 8.39e-07 wmax = 8.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.06983901824397+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.11071507046776
+ k2 = {-0.221261446175075+sky130_fd_pr__pfet_01v8_hvt__k2_diff_54}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.309752008404068
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.250694559258463+sky130_fd_pr__pfet_01v8_hvt__voff_diff_54+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.24943499188874+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.21948113761247+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54}
+ etab = -0.0273684881509353
+ u0 = {0.0028217205352961+sky130_fd_pr__pfet_01v8_hvt__u0_diff_54}
+ ua = {-2.33838595896284e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_54}
+ ub = {2.04285173756036e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_54}
+ uc = 8.58364703942434e-14
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {81709.5428748529+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54}
+ a0 = {1.1332999816516+sky130_fd_pr__pfet_01v8_hvt__a0_diff_54}
+ ags = {1.25000000856918+sky130_fd_pr__pfet_01v8_hvt__ags_diff_54}
+ a1 = 0.0
+ a2 = 0.645206550408959
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_54}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_54}
+ keta = {0.000774133574642732+sky130_fd_pr__pfet_01v8_hvt__keta_diff_54}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.622076876838991+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54}
+ pdiblc1 = 0.167730384011285
+ pdiblc2 = 0.00385905435402245
+ pdiblcb = -0.379687613491591
+ drout = 1.00000015593246
+ pscbe1 = 800000000.056997
+ pscbe2 = 7.37820873129092e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35145700583427
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {2.2929704297289e-10+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54}
+ bgidl = {1000000043.63208+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.536270002860088+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54}
+ kt2 = -0.0962590027256385
+ at = 41259.0011413909
+ ute = -0.0500000411568378
+ ua1 = 7.43579873322196e-10
+ ub1 = -4.72600108632185e-19
+ uc1 = -2.1939001841099e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos
* Model Flag Parameters
+ lmin = 1.79e-07 lmax = 1.81e-07 wmin = 1.679e-06 wmax = 1.681e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07581019562893+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.961428255393082
+ k2 = {-0.162005866831761+sky130_fd_pr__pfet_01v8_hvt__k2_diff_55}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.562303405039308
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.257872947389937+sky130_fd_pr__pfet_01v8_hvt__voff_diff_55+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9870370822327+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55}
+ etab = -0.000625
+ u0 = {0.0037413403490566+sky130_fd_pr__pfet_01v8_hvt__u0_diff_55}
+ ua = {-2.09956058459119e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_55}
+ ub = {1.86166461966667e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_55}
+ uc = -8.324553995283e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {118371.997325472+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55}
+ a0 = {0.758099999261006+sky130_fd_pr__pfet_01v8_hvt__a0_diff_55}
+ ags = {1.24999997272013+sky130_fd_pr__pfet_01v8_hvt__ags_diff_55}
+ a1 = 0.0
+ a2 = 0.662874470440252
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_55}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_55}
+ keta = {-0.0730519999606918+sky130_fd_pr__pfet_01v8_hvt__keta_diff_55}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.734690420259434+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55}
+ pdiblc1 = 0.461536473183962
+ pdiblc2 = 0.00987941513820755
+ pdiblcb = -0.224616327814465
+ drout = 0.684413503600629
+ pscbe1 = 800000000.518868
+ pscbe2 = 9.31998164677673e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.94639467130503
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {3.20550031084906e-10+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55}
+ bgidl = {999999975.393082+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.515879992940252+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55}
+ kt2 = -0.0487919994941038
+ at = 9870.39612421382
+ ute = -0.0199999991650943
+ ua1 = 8.53380055896226e-10
+ ub1 = -4.69150049528303e-19
+ uc1 = -2.62609955581761e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 3.59e-07 wmax = 3.61e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.0751186382512+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.915817576187918
+ k2 = {-0.191354581465138+sky130_fd_pr__pfet_01v8_hvt__k2_diff_56}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.632029034401906
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.252068561266462+sky130_fd_pr__pfet_01v8_hvt__voff_diff_56+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.06838122728761+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.709002668530266+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56}
+ etab = 0.0119734813782515
+ u0 = {0.00388572612584648+sky130_fd_pr__pfet_01v8_hvt__u0_diff_56}
+ ua = {-2.00244775464247e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_56}
+ ub = {1.8126637343077e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_56}
+ uc = -3.29420596540557e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {123538.047249085+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56}
+ a0 = {0.999069843161314+sky130_fd_pr__pfet_01v8_hvt__a0_diff_56}
+ ags = {1.24999999958161+sky130_fd_pr__pfet_01v8_hvt__ags_diff_56}
+ a1 = 0.0
+ a2 = 0.402340703539025
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_56}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_56}
+ keta = {-0.059104614991198+sky130_fd_pr__pfet_01v8_hvt__keta_diff_56}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.626485556768748+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56}
+ pdiblc1 = 0.156960184691247
+ pdiblc2 = 0.00484688249504905
+ pdiblcb = -0.816101282025912
+ drout = 0.999999999574636
+ pscbe1 = 813825374.586324
+ pscbe2 = 9.67821053778591e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.66184153982975
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56}
+ bgidl = {1000000000.29118+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.486150550825388+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56}
+ kt2 = -0.0168844133026869
+ at = 23782.3869663337
+ ute = -0.163199999725863
+ ua1 = 9.15790453404767e-10
+ ub1 = -6.16621741789699e-19
+ uc1 = -1.12531129150376e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 5.39e-07 wmax = 5.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07193945626403+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.04559183372851
+ k2 = {-0.215394224823221+sky130_fd_pr__pfet_01v8_hvt__k2_diff_57}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.296842320875032
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.295820509983861+sky130_fd_pr__pfet_01v8_hvt__voff_diff_57+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.37678785711657+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.203241924319623+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57}
+ etab = -0.0171212205536331
+ u0 = {0.00323243409794057+sky130_fd_pr__pfet_01v8_hvt__u0_diff_57}
+ ua = {-2.18318076500906e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_57}
+ ub = {1.98261706093836e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_57}
+ uc = -1.1166432829987e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {95226.0713945394+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57}
+ a0 = {1.01271311354065+sky130_fd_pr__pfet_01v8_hvt__a0_diff_57}
+ ags = {1.24999999958161+sky130_fd_pr__pfet_01v8_hvt__ags_diff_57}
+ a1 = 0.0
+ a2 = 0.937616983056422
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_57}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_57}
+ keta = {0.0375836653953772+sky130_fd_pr__pfet_01v8_hvt__keta_diff_57}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.622064900782435+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57}
+ pdiblc1 = 0.171475423595225
+ pdiblc2 = 0.00221173256568527
+ pdiblcb = -0.100536440190325
+ drout = 0.999999999572752
+ pscbe1 = 781896315.787039
+ pscbe2 = 9.20129159085351e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.01546307141611
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57}
+ bgidl = {1000000000.29118+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.569263924940705+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57}
+ kt2 = -0.0905365684029605
+ at = 54653.3062207582
+ ute = -0.163199999620793
+ ua1 = 7.49513926681154e-10
+ ub1 = -6.46339460623668e-19
+ uc1 = -4.38452014066302e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 6.29e-07 wmax = 6.31e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07104001525555+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.06962463166075
+ k2 = {-0.211623873447702+sky130_fd_pr__pfet_01v8_hvt__k2_diff_58}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.419583614144431
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.29507245959929+sky130_fd_pr__pfet_01v8_hvt__voff_diff_58+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.23204351258518+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.460564927265331+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58}
+ etab = -0.00252312162912138
+ u0 = {0.00270856257428232+sky130_fd_pr__pfet_01v8_hvt__u0_diff_58}
+ ua = {-2.35623809165088e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_58}
+ ub = {2.04416033113035e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_58}
+ uc = -1.20430539022406e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {85296.9435202141+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58}
+ a0 = {0.890270208902574+sky130_fd_pr__pfet_01v8_hvt__a0_diff_58}
+ ags = {1.25000000001081+sky130_fd_pr__pfet_01v8_hvt__ags_diff_58}
+ a1 = 0.0
+ a2 = 0.768782773323293
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_58}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_58}
+ keta = {-0.00738082267404039+sky130_fd_pr__pfet_01v8_hvt__keta_diff_58}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.620881601802915+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58}
+ pdiblc1 = 0.337392702882825
+ pdiblc2 = 0.00132216097657461
+ pdiblcb = -1.03630654165047
+ drout = 0.999999999645444
+ pscbe1 = 798141699.766914
+ pscbe2 = 5.54371049699427e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.31903127511159
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58}
+ bgidl = {1000000000.27512+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.585293605067905+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58}
+ kt2 = -0.0548785185501603
+ at = 21898.9416489813
+ ute = -0.452342938291501
+ ua1 = 3.87989740344634e-10
+ ub1 = -1.65392727017805e-19
+ uc1 = -3.04688147574841e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 6.99e-07 wmax = 7.01e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07055203747247+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.08580882942068
+ k2 = {-0.214793482817612+sky130_fd_pr__pfet_01v8_hvt__k2_diff_59}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.389054614996031
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.278865636416663+sky130_fd_pr__pfet_01v8_hvt__voff_diff_59+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.59179008241638+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.392167002521586+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59}
+ etab = -0.0104414730939175
+ u0 = {0.00271533057175788+sky130_fd_pr__pfet_01v8_hvt__u0_diff_59}
+ ua = {-2.36115028548009e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_59}
+ ub = {2.04747266512321e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_59}
+ uc = -8.47970537223393e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {83391.0155162216+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59}
+ a0 = {0.969773722807888+sky130_fd_pr__pfet_01v8_hvt__a0_diff_59}
+ ags = {1.25000000001081+sky130_fd_pr__pfet_01v8_hvt__ags_diff_59}
+ a1 = 0.0
+ a2 = 0.711267731601041
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_59}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_59}
+ keta = {-0.0077351739167264+sky130_fd_pr__pfet_01v8_hvt__keta_diff_59}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.621243899946381+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59}
+ pdiblc1 = 0.287320383025818
+ pdiblc2 = 0.00218534505453089
+ pdiblcb = -0.864434997791972
+ drout = 0.999999999569002
+ pscbe1 = 799999999.981033
+ pscbe2 = 5.95874362758602e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3530459991552
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59}
+ bgidl = {1000000000.27513+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.568455637988552+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59}
+ kt2 = -0.0672312825069631
+ at = 26590.3412304301
+ ute = -0.326565404147138
+ ua1 = 4.92325198112386e-10
+ ub1 = -2.43604483811876e-19
+ uc1 = -2.66385372292091e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 7.49e-07 wmax = 7.51e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07026603980288+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.09579867425115
+ k2 = {-0.217387760765392+sky130_fd_pr__pfet_01v8_hvt__k2_diff_60}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.357246668535634
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.267566285842438+sky130_fd_pr__pfet_01v8_hvt__voff_diff_60+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.85556990654462+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.322903101140967+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60}
+ etab = -0.0172308393417141
+ u0 = {0.00275800311393476+sky130_fd_pr__pfet_01v8_hvt__u0_diff_60}
+ ua = {-2.35201958584296e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_60}
+ ub = {2.04561928756625e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_60}
+ uc = -5.04408775493168e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {82716.6038226786+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60}
+ a0 = {1.03536371655589+sky130_fd_pr__pfet_01v8_hvt__a0_diff_60}
+ ags = {1.25000000001081+sky130_fd_pr__pfet_01v8_hvt__ags_diff_60}
+ a1 = 0.0
+ a2 = 0.684770751621682
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_60}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_60}
+ keta = {-0.00432212074264378+sky130_fd_pr__pfet_01v8_hvt__keta_diff_60}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.62157801025884+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60}
+ pdiblc1 = 0.239353130407191
+ pdiblc2 = 0.00285666674423421
+ pdiblcb = -0.670003950087693
+ drout = 0.999999999569002
+ pscbe1 = 799999999.981033
+ pscbe2 = 6.52808779145287e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35240881580645
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60}
+ bgidl = {1000000000.27513+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.555546056520191+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60}
+ kt2 = -0.0788742297123681
+ at = 32473.9047482058
+ ute = -0.21563569030694
+ ua1 = 5.93102890797911e-10
+ ub1 = -3.3545403082025e-19
+ uc1 = -2.47535642267383e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 7.89e-07 wmax = 7.91e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07006394020185+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.10285797531987
+ k2 = {-0.219221001361228+sky130_fd_pr__pfet_01v8_hvt__k2_diff_61}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.334769655703878
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.259581625526074+sky130_fd_pr__pfet_01v8_hvt__voff_diff_61+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.0419693177443+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.273957923178976+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61}
+ etab = -0.0220285295183251
+ u0 = {0.00278815756855406+sky130_fd_pr__pfet_01v8_hvt__u0_diff_61}
+ ua = {-2.34556739776593e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_61}
+ ub = {2.04430960254203e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_61}
+ uc = -2.61631640020886e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {82240.0323373573+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61}
+ a0 = {1.08171273606723+sky130_fd_pr__pfet_01v8_hvt__a0_diff_61}
+ ags = {1.25000000001081+sky130_fd_pr__pfet_01v8_hvt__ags_diff_61}
+ a1 = 0.0
+ a2 = 0.666046721142683
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_61}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_61}
+ keta = {-0.00191029450026639+sky130_fd_pr__pfet_01v8_hvt__keta_diff_61}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.621814108549238+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61}
+ pdiblc1 = 0.205457180728222
+ pdiblc2 = 0.00333105468538863
+ pdiblcb = -0.53260969360584
+ drout = 0.999999999569001
+ pscbe1 = 799999999.981033
+ pscbe2 = 6.93041354652335e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35195855164609
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61}
+ bgidl = {1000000000.27513+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.546423530214438+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61}
+ kt2 = -0.0871016918046216
+ at = 36631.5114912298
+ ute = -0.137247460984637
+ ua1 = 6.64317217521819e-10
+ ub1 = -4.00359303761043e-19
+ uc1 = -2.34215523530136e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 8.19e-07 wmax = 8.21e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.06992560723304+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.1076899199134
+ k2 = {-0.220475816377538+sky130_fd_pr__pfet_01v8_hvt__k2_diff_62}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.319384608434502
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.254116291795267+sky130_fd_pr__pfet_01v8_hvt__voff_diff_62+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.16955583352185+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.24045596799526+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62}
+ etab = -0.0253124485472229
+ u0 = {0.00280879766486815+sky130_fd_pr__pfet_01v8_hvt__u0_diff_62}
+ ua = {-2.34115100937397e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_62}
+ ub = {2.04341315041308e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_62}
+ uc = -9.54557458696919e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {81913.8290787754+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62}
+ a0 = {1.11343767484841+sky130_fd_pr__pfet_01v8_hvt__a0_diff_62}
+ ags = {1.25000000001081+sky130_fd_pr__pfet_01v8_hvt__ags_diff_62}
+ a1 = 0.0
+ a2 = 0.653230512149571
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_62}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_62}
+ keta = {-0.000259449656147479+sky130_fd_pr__pfet_01v8_hvt__keta_diff_62}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.621975712913002+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62}
+ pdiblc1 = 0.182256108950811
+ pdiblc2 = 0.00365576335345378
+ pdiblcb = -0.438566185852545
+ drout = 0.999999999569001
+ pscbe1 = 799999999.981033
+ pscbe2 = 7.20579714868519e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35165035520367
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62}
+ bgidl = {1000000000.27513+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.540179350906419+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62}
+ kt2 = -0.0927332182954322
+ at = 39477.3067375863
+ ute = -0.0835923502048591
+ ua1 = 7.1306194134723e-10
+ ub1 = -4.44785611638355e-19
+ uc1 = -2.25098179604581e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos
* Model Flag Parameters
+ lmin = 1.79e-07 lmax = 1.81e-07 wmin = 8.19e-07 wmax = 8.21e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.06992562425025+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.10768988287566
+ k2 = {-0.220475829959917+sky130_fd_pr__pfet_01v8_hvt__k2_diff_63}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.319384288778231
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.254116290690764+sky130_fd_pr__pfet_01v8_hvt__voff_diff_63+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.16955569641286+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.240456012141059+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63}
+ etab = -0.0253124918524043
+ u0 = {0.00280879816148047+sky130_fd_pr__pfet_01v8_hvt__u0_diff_63}
+ ua = {-2.34115097548295e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_63}
+ ub = {2.04341299867443e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_63}
+ uc = -9.54556263358326e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {81913.7762607886+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63}
+ a0 = {1.11343767246333+sky130_fd_pr__pfet_01v8_hvt__a0_diff_63}
+ ags = {1.25000000883084+sky130_fd_pr__pfet_01v8_hvt__ags_diff_63}
+ a1 = 0.0
+ a2 = 0.653230512297813
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_63}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_63}
+ keta = {-0.000259427474019525+sky130_fd_pr__pfet_01v8_hvt__keta_diff_63}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.621975700968687+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63}
+ pdiblc1 = 0.182256099041279
+ pdiblc2 = 0.00365576108529427
+ pdiblcb = -0.438566290778736
+ drout = 1.00000014412332
+ pscbe1 = 800000000.092367
+ pscbe2 = 7.20579676912272e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.35164997919705
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63}
+ bgidl = {1000000043.76336+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.540179356912575+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63}
+ kt2 = -0.0927332236807995
+ at = 39477.3084346575
+ ute = -0.0835923913034282
+ ua1 = 7.13061837954044e-10
+ ub1 = -4.44785720876955e-19
+ uc1 = -2.25098194407179e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos
* Model Flag Parameters
+ lmin = 2.49e-07 lmax = 2.51e-07 wmin = 8.19e-07 wmax = 8.21e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.05072276049759+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.577863902712096
+ k2 = {-0.0179469684948697+sky130_fd_pr__pfet_01v8_hvt__k2_diff_64}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.784590850821159
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.222875737669666+sky130_fd_pr__pfet_01v8_hvt__voff_diff_64+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.41661831253614+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.490000000534678+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64}
+ etab = -7.18045260867479e-5
+ u0 = {0.00574001096693589+sky130_fd_pr__pfet_01v8_hvt__u0_diff_64}
+ ua = {-1.32599936581963e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_64}
+ ub = {1.3166834291246e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_64}
+ uc = -9.89799750999406e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {96750.2832616657+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64}
+ a0 = {0.615122486656536+sky130_fd_pr__pfet_01v8_hvt__a0_diff_64}
+ ags = {1.50607608496406+sky130_fd_pr__pfet_01v8_hvt__ags_diff_64}
+ a1 = 0.0
+ a2 = 0.796021941247706
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_64}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_64}
+ keta = {-0.0317026683516117+sky130_fd_pr__pfet_01v8_hvt__keta_diff_64}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.637201200109745+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64}
+ pdiblc1 = 0.404629799819182
+ pdiblc2 = 0.00857651181139204
+ pdiblcb = -0.288019851903862
+ drout = 0.528681191381859
+ pscbe1 = 799973295.56758
+ pscbe2 = 8.84471866309014e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.90994629846007
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64}
+ bgidl = {1240180091.56982+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075560999735681*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.47010003888781e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.522777693066561+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64}
+ kt2 = -0.0528131862121549
+ at = 67887.696205111
+ ute = -0.83458849565544
+ ua1 = 2.95036202917305e-10
+ ub1 = -1.69321451147667e-19
+ uc1 = -9.78860164868713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos
* Model Flag Parameters
+ lmin = 4.99e-07 lmax = 5.01e-07 wmin = 8.19e-07 wmax = 8.21e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-1.176e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.05257645277475+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.509746853558371
+ k2 = {0.0010565381342913+sky130_fd_pr__pfet_01v8_hvt__k2_diff_65}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.319727369402999
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.207851692258142+sky130_fd_pr__pfet_01v8_hvt__voff_diff_65+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.07922336976018+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.452641007151395+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65}
+ etab = -0.000654076810703508
+ u0 = {0.00682669236101063+sky130_fd_pr__pfet_01v8_hvt__u0_diff_65}
+ ua = {-1.20060863280976e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_65}
+ ub = {1.23616934688699e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_65}
+ uc = -3.11715075302948e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {98242.5308183485+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65}
+ a0 = {0.747334484184591+sky130_fd_pr__pfet_01v8_hvt__a0_diff_65}
+ ags = {1.24999999994093+sky130_fd_pr__pfet_01v8_hvt__ags_diff_65}
+ a1 = 0.0
+ a2 = 0.951482129181008
+ b0 = {8.77074029519858e-17+sky130_fd_pr__pfet_01v8_hvt__b0_diff_65}
+ b1 = {3.64639825577157e-20+sky130_fd_pr__pfet_01v8_hvt__b1_diff_65}
+ keta = {-0.0381687151274896+sky130_fd_pr__pfet_01v8_hvt__keta_diff_65}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.0592215633585798+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65}
+ pdiblc1 = 0.0155649705144554
+ pdiblc2 = 9.9333572416857e-5
+ pdiblcb = -0.0354604781743123
+ drout = 0.962160634824741
+ pscbe1 = 748693433.4003
+ pscbe2 = 1.4666228889085e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.72758012904933
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65}
+ bgidl = {1000000000.0+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-2.56e-09+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.533868339386531+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65}
+ kt2 = -0.034749082504185
+ at = 38573.0516436388
+ ute = -0.201655304750119
+ ua1 = 2.4966480698116e-9
+ ub1 = -2.31670144462701e-18
+ uc1 = -1.85406901254478e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 8.59e-07 wmax = 8.61e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07104381577694+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.10594770014062
+ k2 = {-0.219965620603534+sky130_fd_pr__pfet_01v8_hvt__k2_diff_66}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.308703572208419
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.257630636013059+sky130_fd_pr__pfet_01v8_hvt__voff_diff_66+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.09352853651824+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.216916404856265+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66}
+ etab = -0.025065060370094
+ u0 = {0.0029364922909248+sky130_fd_pr__pfet_01v8_hvt__u0_diff_66}
+ ua = {-2.2922101231441e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_66}
+ ub = {1.99787255718905e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_66}
+ uc = 7.56985290191209e-14
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {81250.6743978597+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66}
+ a0 = {1.10173536063403+sky130_fd_pr__pfet_01v8_hvt__a0_diff_66}
+ ags = {1.25000000032035+sky130_fd_pr__pfet_01v8_hvt__ags_diff_66}
+ a1 = 0.0
+ a2 = 0.668724680856823
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_66}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_66}
+ keta = {0.000585058556570317+sky130_fd_pr__pfet_01v8_hvt__keta_diff_66}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.622098795779318+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66}
+ pdiblc1 = 0.165599715192776
+ pdiblc2 = 0.00370966311736148
+ pdiblcb = -0.373536489052468
+ drout = 0.999999994584648
+ pscbe1 = 799999999.950522
+ pscbe2 = 7.51810401745175e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.33366985234279
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66}
+ bgidl = {999999999.964758+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.540644055101813+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66}
+ kt2 = -0.0962590000996655
+ at = 38488.7652643574
+ ute = -0.0434389167673217
+ ua1 = 7.43579997969786e-10
+ ub1 = -4.7259999135388e-19
+ uc1 = -2.19389998907211e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos
* Model Flag Parameters
+ lmin = 1.49e-07 lmax = 1.51e-07 wmin = 9.39e-07 wmax = 9.41e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.23e-09*sky130_fd_pr__pfet_01v8_hvt__toxe_mult+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*sky130_fd_pr__pfet_01v8_hvt__toxe_mult*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = {1.0*sky130_fd_pr__pfet_01v8_hvt__rshp_mult}
+ rshg = 0.1
* Basic Model Parameters
+ wint = {9.364e-09+sky130_fd_pr__pfet_01v8_hvt__wint_diff}
+ lint = {-2.026e-08+sky130_fd_pr__pfet_01v8_hvt__lint_diff}
+ vth0 = {-1.07533996982605+sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 1.08894802372141
+ k2 = {-0.215345000473891+sky130_fd_pr__pfet_01v8_hvt__k2_diff_67}
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.304963807285077
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.282363418797658+sky130_fd_pr__pfet_01v8_hvt__voff_diff_67+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.53759417857265+sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = {0.207771195728855+sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67}
+ etab = -0.0168516215301728
+ u0 = {0.00334574934342391+sky130_fd_pr__pfet_01v8_hvt__u0_diff_67}
+ ua = {-2.12755536041125e-09+sky130_fd_pr__pfet_01v8_hvt__ua_diff_67}
+ ub = {1.83748442782511e-18+sky130_fd_pr__pfet_01v8_hvt__ub_diff_67}
+ uc = 3.95528374555728e-14
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = {79614.2284598555+sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67}
+ a0 = {0.989181612672348+sky130_fd_pr__pfet_01v8_hvt__a0_diff_67}
+ ags = {1.25000000032035+sky130_fd_pr__pfet_01v8_hvt__ags_diff_67}
+ a1 = 0.0
+ a2 = 0.752586056400402
+ b0 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b0_diff_67}
+ b1 = {0.0+sky130_fd_pr__pfet_01v8_hvt__b1_diff_67}
+ keta = {-8.906293497013e-05+sky130_fd_pr__pfet_01v8_hvt__keta_diff_67}
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = {0.622176905948925+sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67}
+ pdiblc1 = 0.158002074710554
+ pdiblc2 = 0.00317695286612851
+ pdiblcb = -0.351603091257726
+ drout = 0.999999995175411
+ pscbe1 = 799999999.950522
+ pscbe2 = 8.01694390444676e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = {0.0+sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67}
+ pditsl = 0.0
+ pditsd = {0.0+sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67}
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = {531.92+sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67}
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.27024270366315
* Gidl Induced Drain Leakage Model Parameters
+ agidl = {0.0+sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67}
+ bgidl = {999999999.964757+sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67}
+ cgidl = {300.0+sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67}
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = {-1.106e-08+sky130_fd_pr__pfet_01v8_hvt__dlc_diff+sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak}
+ dwc = {0.0+sky130_fd_pr__pfet_01v8_hvt__dwc_diff}
+ xpart = 0.0
+ cgso = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgdo = {6.0e-11*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgbo = 0.0
+ cgdl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ cgsl = {7.6e-12*sky130_fd_pr__pfet_01v8_hvt__overlap_mult}
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = {0.00075561*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult}
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = {9.2435e-11*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = {2.4701e-10*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult}
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = {-0.556241137832508+sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67}
+ kt2 = -0.096259000063518
+ at = 28610.6128567872
+ ute = -0.0200432924793255
+ ua1 = 7.43579998498136e-10
+ ub1 = -4.72599991749167e-19
+ uc1 = -2.19389998945569e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = {0.0+sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67}
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
.ends sky130_fd_pr__pfet_01v8_hvt
* Well Proximity Effect Parameters
