* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./models_resistors.spice created from ./models.spice
*
**********************************
******************************************************************
******************************************************************
***************************************************************************
**
**   Interconnect, parasitic and misc resistors
**
***************************************************************************


**  resistance temperature coeff
**All the way up to M1 is the same between these technologies, so all those files are the same here

.param   tc1rsn=  1.422E-03
.param   tc2rsn=  6.569e-7
.param   tc1rsp=   1.259e-3
.param   tc2rsp=   2.204e-6 
.param   tc1rsn_h=  1.405E-03
.param   tc2rsn_h=  4.233e-7
.param   tc1rsp_h=   1.369e-3
.param   tc2rsp_h=   1.476e-6
.param   tc1rsnw=  1.483e-3
.param   tc2rsnw=  7.824e-6
.param   tc1rsgpw= 8.100e-04
.param   tc2rsgpw= 7.840e-7
.param   tc1rsgpu= 8.916e-4
.param   tc2rsgpu= 8.443e-7

.param   tc1rl1=   6.045e-4
.param   tc2rl1=  -3.693e-7
.param   tc1sky130_fd_pr__res_generic_m1=   3.179e-3
.param   tc2sky130_fd_pr__res_generic_m1=   3.094e-7
.param   tc1sky130_fd_pr__res_generic_m2=   3.161e-3
.param   tc2sky130_fd_pr__res_generic_m2=  -7.272e-7
.param   tc1sky130_fd_pr__res_generic_m3=   3.424e-3
.param   tc2sky130_fd_pr__res_generic_m3=  -7.739e-7
.param   tc1sky130_fd_pr__res_generic_m4=   3.424e-3
.param   tc2sky130_fd_pr__res_generic_m4=  -7.739e-7
.param   tc1sky130_fd_pr__res_generic_m5=   3.500e-3
.param   tc2sky130_fd_pr__res_generic_m5=  -7.500e-7
.param   tc1rrdl=  3.930e-3
.param   tc2rrdl=  0.0

.param   tc1rcn=   2.254e-4
.param   tc2rcn=  -1.038e-6
.param   tc1rcp=   5.250e-4
.param   tc2rcp=   3.544e-6
.param   tc1rcgp=  1.249e-3
.param   tc2rcgp= -6.647e-6
.param   tc1rcl1=  1.067e-3
.param   tc2rcl1= -5.324e-6
.param   tc1rvia=  1.081e-3
.param   tc2rvia= -1.903e-7
.param   tc1rvia2= 2.366e-3
.param   tc2rvia2=-1.025e-5
.param   tc1rvia3= 2.366e-3
.param   tc2rvia3=-1.025e-5
.param   tc1rvia4= 1.77e-03
.param   tc2rvia4= -1.60e-07
.param   tc1rrdlcon=  3.930e-3
.param   tc2rrdlcon=  0.0

.param   tc1sky130_fd_pr__res_generic_pobody= 0.514e-3
.param   tc2sky130_fd_pr__res_generic_pobody= 0.122e-5
.param   tc1sky130_fd_pr__res_generic_poend=  0.0
.param   tc2sky130_fd_pr__res_generic_poend=  0.0

* +     sw_tc1sky130_fd_pr__res_generic_m3     = 3.424e-3   sw_tc2sky130_fd_pr__res_generic_m3   = -7.739e-7
* +     sw_tc1sky130_fd_pr__res_generic_m4     = 3.424e-3   sw_tc2sky130_fd_pr__res_generic_m4   = -7.739e-7
* +     sw_tc1rvia3   = 2.366e-3   sw_tc2rvia3 = -1.025e-5
* +     sw_tc1rvia4   = 1.77e-03   sw_tc2rvia4 = -1.60e-07

***************************************
* differences between the electrical  *
*      and scaled drawn widths        *
***************************************
.param
+ nfom_dw = 0.017u
+ pfom_dw = 0.004u
+ poly_dw = -0.056u
+ li_dw =  0.017u
+ m1_dw = -0.039u
+ m2_dw = -0.039u
+ m3_dw = -0.025u
+ m4_dw = -0.025u
+ m5_dw = -0.09u
+ rdl_dw = 0.0u


********************************************************************
*          model for interconnect resistance       *
********************************************************************

.model rndiff r tc1 = {tc1rsn} tc2 = {tc2rsn} rsh = {sw_rdn} dw = {"-sw_activecd-nfom_dw/2"} tref = 30
.model rpdiff r tc1 = {tc1rsp} tc2 = {tc2rsp} rsh = {sw_rdp} dw = {"-sw_activecd-pfom_dw/2"} tref = 30
.model rndiff_v5 r tc1 = {tc1rsn_h} tc2 = {tc2rsn_h} rsh = {sw_rdn*0.95} dw = {"-sw_activecd-nfom_dw/2"} tref = 30
.model rpdiff_v5 r tc1 = {tc1rsp_h} tc2 = {tc2rsp_h} rsh = {sw_rdp*0.97} dw = {"-sw_activecd-pfom_dw/2"} tref = 30
.model rnwell r tc1 = {tc1rsnw} tc2 = {tc2rsnw} rsh = {sw_rnw} dw = {"-sw_activecd/2"} tref = 30
.model sky130_fd_pr__res_generic_l1 r tc1 = {tc1rl1} tc2 = {tc2rl1} rsh = {sw_rl1} dw = {"-sw_rl1_dw/2-li_dw/2"} tref = 30
.model sky130_fd_pr__res_generic_m1 r tc1 = {tc1sky130_fd_pr__res_generic_m1} tc2 = {tc2sky130_fd_pr__res_generic_m1} rsh = {sw_sky130_fd_pr__res_generic_m1_rs} dw = {"-sw_m1_dw/2-m1_dw/2"} tref = 30
.model sky130_fd_pr__res_generic_m2 r tc1 = {tc1sky130_fd_pr__res_generic_m2} tc2 = {tc2sky130_fd_pr__res_generic_m2} rsh = {sw_sky130_fd_pr__res_generic_m2_rs} dw = {"-sw_m2_dw/2-m2_dw/2"} tref = 30
.model sky130_fd_pr__res_generic_m3 r tc1 = {tc1sky130_fd_pr__res_generic_m3} tc2 = {tc2sky130_fd_pr__res_generic_m3} rsh = {sw_sky130_fd_pr__res_generic_m3_rs} dw = {"-sw_m3_dw/2-m3_dw/2"} tref = 30
.model sky130_fd_pr__res_generic_m4 r tc1 = {tc1sky130_fd_pr__res_generic_m4} tc2 = {tc2sky130_fd_pr__res_generic_m4} rsh = {sw_sky130_fd_pr__res_generic_m4_rs} dw = {"-sw_m4_dw/2-m4_dw/2"} tref = 30
.model sky130_fd_pr__res_generic_m5 r tc1 = {tc1sky130_fd_pr__res_generic_m5} tc2 = {tc2sky130_fd_pr__res_generic_m5} rsh = {sw_sky130_fd_pr__res_generic_m5_rs} dw = {"-sw_m5_dw/2-m5_dw/2"} tref = 30
.model mrrdl r tc1 = {tc1rrdl} tc2 = {tc2rrdl} rsh = {rrdl} dw = {"-tol_rdl/2-rdl_dw/2"} tref = 25
.model mrcn r tc1 = {tc1rcn} tc2 = {tc2rcn} res = {rcn} tref = 30
.model mrcp r tc1 = {tc1rcp} tc2 = {tc2rcp} res = {rcp} tref = 30
.model mrcp1 r tc1 = {tc1rcgp} tc2 = {tc2rcgp} res = {rcp1} tref = 30
.model mrcl1 r tc1 = {tc1rcl1} tc2 = {tc2rcl1} res = {rcl1} tref = 30
.model mrcvia r tc1 = {tc1rvia} tc2 = {tc2rvia} res = {rcvia} tref = 30
.model mrcvia2 r tc1 = {tc1rvia2} tc2 = {tc2rvia2} res = {rcvia2} tref = 30
.model mrcvia3 r tc1 = {tc1rvia3} tc2 = {tc2rvia3} res = {rcvia3} tref = 30
.model mrcvia4 r tc1 = {tc1rvia4} tc2 = {tc2rvia4} res = {rcvia4} tref = 30
.model mrcrdlcon r tc1 = {tc1rrdlcon} tc2 = {tc2rrdlcon} res = {rcrdlcon} tref = 25

********************************************************************
*          Subcircuit model
********************************************************************

.subckt  sky130_fd_pr__res_generic_nd t1 t2 b mult=1
+ w=1 l=1

r0 t1 t2 rndiff w = {w} l = {l}
xd0 b t1 sky130_fd_pr__diode_pw2nd_05v5 area = 'w*l*0.5' perim = 'w+l'
xd1 b t2 sky130_fd_pr__diode_pw2nd_05v5 area = 'w*l*0.5' perim = 'w+l'

.ends sky130_fd_pr__res_generic_nd

.subckt  sky130_fd_pr__res_generic_pd t1 t2 b mult=1
+ w=1 l=1

r0 t1 t2 rpdiff w = {w} l = {l}
xd0 t1 b sky130_fd_pr__model__parasitic__diode_pd2nw area = 'w*l*0.5' perim = 'w+l'
xd1 t2 b sky130_fd_pr__model__parasitic__diode_pd2nw area = 'w*l*0.5' perim = 'w+l'

.ends sky130_fd_pr__res_generic_pd
******************************************************************
******************************************************************
* *************************** 2K Ohm/sq Poly Resistors ************************
* 2021/03/04  UZMN (Usman Suriono)
*      Why  : New 2K Ohm/sq Poly resistor model
*      What : Data taken from lot 4936073 wafer 11 with 1.4K ohm/sq
*             The model will be updated with 2K ohm/sq silicon in the future.

.subckt  sky130_fd_pr__res_xhigh_po r0 r1 sub mult=1
+ w=1 l=1
* Effective length and width
+ 
.param  leff = {l-0.0592}
+ weff = {w-0.056+2*sw_polycd}
* Resistor voltco fitting parameters
+ bp2 = -0.1228
+ bq2 = 1.304
+ bp22 = -0.2874
+ bp23 = 0.5252
* Substrate voltco fitting parameters
+ sub1 = 1.2 ;  y-axis offset
+ sub2 = 41.26e-3 ;  top-bottom scale
+ sub3 = 8.697e-3 ;  slope of tanh
+ sub4 = 24 ;  half of the plateau voltage (12V)
+ sub5 = 39.86 ;  offset voltage of tanh function
* Resistor head and body scalable equation
+ rhead0 = {188.2/(weff-0.0672*max(0.69-w,0)+1.41)}
+ rbody0 = {sw_sky130_fd_pr__res_xhigh_po_rs*leff/(weff-0.0672*max(0.69-w,0))} ;  the last term for w<0.69 current crowding
* Equations with variation
+ Efac = {1/leff*(1+bp22/w+bp23*min(0.2,leff-0.5)*log(leff/w))}
+ rhead = {rhead0*sw_poly_head_res*(1+sw_mm_sky130_fd_pr__res_generic_po_head*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*mult))}
+ rbody = {rbody0*(1+sw_mm_sky130_fd_pr__res_xhigh_po*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*l*mult))}

rend1 r0 t1 reshead r = {rhead}
rend2 t2 r1 reshead r = {rhead}
xc0 r0 sub sky130_fd_pr__model__parasitic__cap_p2ps w = {weff} l = {l+2.08} m = 0.5
xc1 r1 sub sky130_fd_pr__model__parasitic__cap_p2ps w = {weff} l = {l+2.08} m = 0.5

rbody t1 t2 resbody r = {rbody*(1-bp2+bp2*sqrt(1+(bq2*abs(v(t1,t2))*Efac)**2))*
+ (sub1+sub2*tanh(sub3*(min(v(sub,r1)+v(sub,r1),sub4)+sub5))) / (sub1+sub2*tanh(sub3*sub5)) }


.model resbody r tc1 = {-1.47e-3-5e-7*sw_sky130_fd_pr__res_xhigh_po_rs} tc2 = 2.7e-6 tnom = 25

.model reshead r tc1 = -4.3e-4 tc2 = -1.3e-5 tnom = 25

.ends sky130_fd_pr__res_xhigh_po

******************************************************************
******************************************************************
* *************************** 300 Ohm/sq Scalable Poly Resistors ************************
* 2021/09/03  UZMN (Usman Suriono)
*      Why  : Missing temperature coefficients
*      What : Add temperature coefficients from the original model.
* 2021/03/04  UZMN (Usman Suriono)
*      Why  : New scalable 300 Ohm/sq Poly resistor model
*      What : Converted from discrete model


.subckt  sky130_fd_pr__res_high_po r0 r1 b mult=1
+ w=1 l=1

* parameter values:
+ 
.param  rbody_dw = {-0.001+sw_polycd*2e6}
+ rhead_ps = 345.8312
+ num_con_row = {max(floor(0.5+(w-0.33)/0.36),1)}
* resistance. The max() for exception due to exception spacing when w<0.69
+ weff = {w+rbody_dw-0.0672*max(0.69-w,0)+2*sw_polycd}
+ leff = {l+0.247}

rhead r0 rb rhead_model w = {weff+0.1558} l = 1
rbody rb r1 rbody_model w = {weff} l = {leff}

xc0 r0 b sky130_fd_pr__model__parasitic__cap_p2ps w = {weff} l = {l+2.08} m = 0.5
xc1 r1 b sky130_fd_pr__model__parasitic__cap_p2ps w = {weff} l = {l+2.08} m = 0.5

.model rhead_model r 
+ rsh = {rhead_ps*sw_poly_head_res*(1+sw_mm_sky130_fd_pr__res_generic_po_head*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*mult))}

.model rbody_model r 
+ rsh = {sw_sky130_fd_pr__res_high_po_rs*(1+sw_mm_sky130_fd_pr__res_high_po*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*l*mult))}
+ tc1 = {tc1sky130_fd_pr__res_generic_pobody} tc2 = {tc2sky130_fd_pr__res_generic_pobody} tnom = 30

*   Voltage coefficient models to be verified in the future
*   model rhead_model r2 sw_et=no isnoisy=no
*        + rsh = rhead_ps * sw_poly_head_res * (1+rend_match)
*        + p2  = -80.87e-3 / cosh(6.34e-3* weff*weff ) * (1-exp(-1.554 / leff))
*        + q2  = 10.13 / cosh(0.0898*weff*weff)
*        + tc1=-4.3e-4    tc2=12e-6   tnom=30

*   model rbody_model r2 sw_et=no isnoisy=no
*        + rsh= sw_sky130_fd_pr__res_high_po_rs  * (1 + res_match)
*        + p2 = (w > 0.6)? 130.8e3*(1-exp(-1.818e-3*leff/weff))-867.4/weff+2236*weff/leff : 300*(1-exp(-0.1124*leff/weff))+304.8*weff/leff
*        + q2 = (w > 0.6)? 6.11*(1-exp(-852.8e-6*leff/weff))+1.375e-3*weff : 0.5*0.3155 *(1-exp(-0.05518*leff/weff))+1.19E-05*weff
*        + p3 = (w > 0.6)?  380.3 * weff / leff : 0
*        + q3 = (w > 0.6)? 42.62e-3 * weff / leff : 0


.ends sky130_fd_pr__res_high_po
******************************************************************
******************************************************************
* *************************** 48 Ohm/sq Scalable Poly Resistors ************************
* 2021/03/04  UZMN (Usman Suriono)
*      What : Copied from "sky130_fd_pr__res_generic_po" model
*             Added matching.


.subckt  sky130_fd_pr__res_generic_po r0 r1 mult=1
+ 
.param  w = 1 l = 0 r = 0 tc1 = {tc1rsgpu} tc2 = {tc2rsgpu}
+ r_tot = {sw_rp1*l/(w-1e6*(sw_polycd*4-poly_dw))+r}

Rsky130_fd_pr__res_generic_po r0 r1 r = {r_tot*(1+sw_mm_sky130_fd_pr__res_generic_po*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*l*mult))}
+ tc1 = {tc1} tc2 = {tc2}


.ends sky130_fd_pr__res_generic_po

******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/03/04  UZMN (Usman Suriono)
*      What : Pwell resistor model copied from model
*             Add pwell to Deep Nwell parasitic diode
*             The voltage coefficient from Nwell bias is not modeled yet.
*             Add matching.

.subckt  sky130_fd_pr__res_iso_pw r0 r1 b mult=1
+ 
.param  l = -1 w = 2.65
+ dl = 0.52
+ av = 0.0133
+ bv = 0.0302
+ tref = 30.0
+ vvt = 3.531e-3
+ ut = 7.238e-6
+ rtot = {sw_pw_rs*(1+sw_mm_sky130_fd_pr__res_iso_pw*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(w*l*mult))}

xdnw1 r0 b sky130_fd_pr__model__parasitic__diode_pw2dn area = {(l+dl)*w*0.5} perim = {(l+dl+w)}
xdnw2 r1 b sky130_fd_pr__model__parasitic__diode_pw2dn area = {(l+dl)*w*0.5} perim = {(l+dl+w)}
Rsky130_fd_pr__res_iso_pw r0 r1
+ r = {rtot*sw_pw_rs_mc*((l+dl)/w)*(1-av*(max(v(r0),v(r1))-min(v(r0),v(r1))))*(1+bv*(v(b)-min(v(r0),v(r1))))*(1+vvt*(temper-tref)+ut*(temper-tref)*(temper-tref))}



.ends sky130_fd_pr__res_iso_pw
