# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__ind_01_04
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__ind_01_04 ;
  ORIGIN  98.30000  8.265000 ;
  SIZE  196.6000 BY  164.9150 ;
  PIN CENTERTAP
    PORT
      LAYER met5 ;
        POLYGON -72.500000  35.175000 -64.615000  35.175000 -64.615000  27.290000 ;
        POLYGON -69.335000 115.980000 -69.335000 112.815000 -72.500000 112.815000 ;
        POLYGON -66.500000  37.655000 -64.500000  35.655000 -66.500000  35.655000 ;
        POLYGON -66.500000 112.635000 -64.200000 112.635000 -66.500000 110.335000 ;
        POLYGON -64.615000  27.290000 -57.655000  27.290000 -57.655000  20.330000 ;
        POLYGON -64.500000  35.655000 -61.780000  32.935000 -64.500000  32.935000 ;
        POLYGON -64.500000  38.505000 -63.650000  38.505000 -63.650000  37.655000 ;
        POLYGON -64.200000 115.485000 -61.350000 115.485000 -64.200000 112.635000 ;
        POLYGON -63.650000  37.655000 -61.650000  37.655000 -61.650000  35.655000 ;
        POLYGON -63.650000 110.335000 -63.650000 109.485000 -64.500000 109.485000 ;
        POLYGON -61.780000  32.935000 -60.340000  31.495000 -61.780000  31.495000 ;
        POLYGON -61.650000  35.655000 -58.930000  35.655000 -58.930000  32.935000 ;
        POLYGON -61.350000 112.635000 -61.350000 110.335000 -63.650000 110.335000 ;
        POLYGON -61.350000 118.335000 -58.500000 118.335000 -61.350000 115.485000 ;
        POLYGON -61.350000 123.965000 -61.350000 115.980000 -69.335000 115.980000 ;
        POLYGON -60.340000  31.495000 -57.985000  29.140000 -60.340000  29.140000 ;
        POLYGON -58.930000  32.935000 -57.490000  32.935000 -57.490000  31.495000 ;
        POLYGON -58.500000  40.985000 -56.500000  38.985000 -58.500000  38.985000 ;
        POLYGON -58.500000 107.535000 -57.970000 107.535000 -58.500000 107.005000 ;
        POLYGON -58.500000 115.485000 -58.500000 112.635000 -61.350000 112.635000 ;
        POLYGON -58.500000 121.115000 -55.720000 121.115000 -58.500000 118.335000 ;
        POLYGON -57.985000  29.140000 -56.135000  27.290000 -57.985000  27.290000 ;
        POLYGON -57.970000 110.335000 -55.170000 110.335000 -57.970000 107.535000 ;
        POLYGON -57.655000  20.330000 -52.820000  20.330000 -52.820000  15.495000 ;
        POLYGON -57.490000  31.495000 -55.135000  31.495000 -55.135000  29.140000 ;
        POLYGON -56.500000  38.985000 -55.170000  37.655000 -56.500000  37.655000 ;
        POLYGON -56.500000  41.820000 -55.665000  41.820000 -55.665000  40.985000 ;
        POLYGON -56.135000  27.290000 -53.300000  24.455000 -56.135000  24.455000 ;
        POLYGON -55.720000 123.965000 -52.870000 123.965000 -55.720000 121.115000 ;
        POLYGON -55.665000  40.985000 -53.665000  40.985000 -53.665000  38.985000 ;
        POLYGON -55.665000 107.005000 -55.665000 106.170000 -56.500000 106.170000 ;
        POLYGON -55.650000 118.335000 -55.650000 115.485000 -58.500000 115.485000 ;
        POLYGON -55.170000  37.655000 -53.170000  35.655000 -55.170000  35.655000 ;
        POLYGON -55.170000 112.170000 -53.335000 112.170000 -55.170000 110.335000 ;
        POLYGON -55.135000  29.140000 -53.285000  29.140000 -53.285000  27.290000 ;
        POLYGON -55.135000 107.535000 -55.135000 107.005000 -55.665000 107.005000 ;
        POLYGON -53.665000  38.985000 -52.335000  38.985000 -52.335000  37.655000 ;
        POLYGON -53.335000 115.005000 -50.500000 115.005000 -53.335000 112.170000 ;
        POLYGON -53.300000  24.455000 -51.530000  22.685000 -53.300000  22.685000 ;
        POLYGON -53.285000  27.290000 -50.450000  27.290000 -50.450000  24.455000 ;
        POLYGON -53.170000  35.655000 -50.450000  32.935000 -53.170000  32.935000 ;
        POLYGON -52.870000 121.115000 -52.870000 118.335000 -55.650000 118.335000 ;
        POLYGON -52.870000 126.815000 -50.020000 126.815000 -52.870000 123.965000 ;
        POLYGON -52.870000 132.445000 -52.870000 123.965000 -61.350000 123.965000 ;
        POLYGON -52.820000  15.495000 -44.820000  15.495000 -44.820000   7.495000 ;
        POLYGON -52.335000  37.655000 -50.335000  37.655000 -50.335000  35.655000 ;
        POLYGON -52.335000 110.335000 -52.335000 107.535000 -55.135000 107.535000 ;
        POLYGON -51.530000  22.685000 -49.175000  20.330000 -51.530000  20.330000 ;
        POLYGON -50.500000  44.300000 -48.500000  42.300000 -50.500000  42.300000 ;
        POLYGON -50.500000 106.170000 -48.020000 106.170000 -50.500000 103.690000 ;
        POLYGON -50.500000 112.170000 -50.500000 110.335000 -52.335000 110.335000 ;
        POLYGON -50.500000 115.980000 -49.525000 115.980000 -50.500000 115.005000 ;
        POLYGON -50.450000  24.455000 -48.680000  24.455000 -48.680000  22.685000 ;
        POLYGON -50.450000  32.935000 -49.010000  31.495000 -50.450000  31.495000 ;
        POLYGON -50.335000  35.655000 -47.615000  35.655000 -47.615000  32.935000 ;
        POLYGON -50.020000 123.965000 -50.020000 121.115000 -52.870000 121.115000 ;
        POLYGON -50.020000 129.595000 -47.240000 129.595000 -50.020000 126.815000 ;
        POLYGON -49.540000 135.775000 -49.540000 132.445000 -52.870000 132.445000 ;
        POLYGON -49.525000 118.815000 -46.690000 118.815000 -49.525000 115.980000 ;
        POLYGON -49.175000  20.330000 -46.340000  17.495000 -49.175000  17.495000 ;
        POLYGON -49.010000  31.495000 -46.655000  29.140000 -49.010000  29.140000 ;
        POLYGON -48.680000  22.685000 -46.325000  22.685000 -46.325000  20.330000 ;
        POLYGON -48.500000  42.300000 -45.695000  39.495000 -48.500000  39.495000 ;
        POLYGON -48.500000  45.140000 -47.660000  45.140000 -47.660000  44.300000 ;
        POLYGON -48.020000 108.850000 -45.340000 108.850000 -48.020000 106.170000 ;
        POLYGON -48.015000 103.335000 -48.015000 102.850000 -48.500000 102.850000 ;
        POLYGON -47.665000 115.005000 -47.665000 112.170000 -50.500000 112.170000 ;
        POLYGON -47.660000  44.300000 -45.660000  44.300000 -45.660000  42.300000 ;
        POLYGON -47.660000 103.690000 -47.660000 103.335000 -48.015000 103.335000 ;
        POLYGON -47.615000  32.935000 -46.175000  32.935000 -46.175000  31.495000 ;
        POLYGON -47.240000 132.445000 -44.390000 132.445000 -47.240000 129.595000 ;
        POLYGON -47.170000 126.815000 -47.170000 123.965000 -50.020000 123.965000 ;
        POLYGON -46.820000 138.495000 -46.820000 135.775000 -49.540000 135.775000 ;
        POLYGON -46.690000 115.980000 -46.690000 115.005000 -47.665000 115.005000 ;
        POLYGON -46.690000 120.650000 -44.855000 120.650000 -46.690000 118.815000 ;
        POLYGON -46.655000  29.140000 -44.805000  27.290000 -46.655000  27.290000 ;
        POLYGON -46.340000  17.495000 -44.340000  15.495000 -46.340000  15.495000 ;
        POLYGON -46.325000  20.330000 -43.490000  20.330000 -43.490000  17.495000 ;
        POLYGON -46.175000  31.495000 -43.820000  31.495000 -43.820000  29.140000 ;
        POLYGON -45.695000  39.495000 -42.855000  36.655000 -45.695000  36.655000 ;
        POLYGON -45.660000  42.300000 -42.855000  42.300000 -42.855000  39.495000 ;
        POLYGON -45.340000 111.690000 -42.500000 111.690000 -45.340000 108.850000 ;
        POLYGON -45.180000 106.170000 -45.180000 103.690000 -47.660000 103.690000 ;
        POLYGON -44.855000 122.495000 -43.010000 122.495000 -44.855000 120.650000 ;
        POLYGON -44.820000   7.495000 -38.820000   7.495000 -38.820000   1.495000 ;
        POLYGON -44.805000  27.290000 -41.970000  24.455000 -44.805000  24.455000 ;
        POLYGON -44.390000 129.595000 -44.390000 126.815000 -47.170000 126.815000 ;
        POLYGON -44.390000 135.295000 -41.540000 135.295000 -44.390000 132.445000 ;
        POLYGON -44.340000  15.495000 -41.490000  12.645000 -44.340000  12.645000 ;
        POLYGON -43.855000 118.815000 -43.855000 115.980000 -46.690000 115.980000 ;
        POLYGON -43.820000  29.140000 -41.970000  29.140000 -41.970000  27.290000 ;
        POLYGON -43.490000  17.495000 -41.490000  17.495000 -41.490000  15.495000 ;
        POLYGON -43.010000 124.495000 -41.010000 124.495000 -43.010000 122.495000 ;
        POLYGON -42.855000  36.655000 -40.505000  34.305000 -42.855000  34.305000 ;
        POLYGON -42.855000  39.495000 -40.015000  39.495000 -40.015000  36.655000 ;
        POLYGON -42.855000 108.495000 -42.855000 106.170000 -45.180000 106.170000 ;
        POLYGON -42.500000  47.620000 -40.500000  45.620000 -42.500000  45.620000 ;
        POLYGON -42.500000 100.495000 -42.375000 100.495000 -42.500000 100.370000 ;
        POLYGON -42.500000 108.850000 -42.500000 108.495000 -42.855000 108.495000 ;
        POLYGON -42.500000 114.495000 -39.695000 114.495000 -42.500000 111.690000 ;
        POLYGON -42.375000 103.335000 -39.535000 103.335000 -42.375000 100.495000 ;
        POLYGON -42.020000 120.650000 -42.020000 118.815000 -43.855000 118.815000 ;
        POLYGON -41.970000  24.455000 -40.200000  22.685000 -41.970000  22.685000 ;
        POLYGON -41.970000  27.290000 -39.135000  27.290000 -39.135000  24.455000 ;
        POLYGON -41.540000 132.445000 -41.540000 129.595000 -44.390000 129.595000 ;
        POLYGON -41.540000 135.775000 -41.060000 135.775000 -41.540000 135.295000 ;
        POLYGON -41.490000  12.645000 -41.190000  12.345000 -41.490000  12.345000 ;
        POLYGON -41.490000  15.495000 -38.640000  15.495000 -38.640000  12.645000 ;
        POLYGON -41.190000  12.345000 -38.340000   9.495000 -41.190000   9.495000 ;
        POLYGON -41.060000 138.495000 -38.340000 138.495000 -41.060000 135.775000 ;
        POLYGON -41.010000 127.295000 -38.210000 127.295000 -41.010000 124.495000 ;
        POLYGON -40.505000  34.305000 -37.695000  31.495000 -40.505000  31.495000 ;
        POLYGON -40.500000  45.620000 -39.180000  44.300000 -40.500000  44.300000 ;
        POLYGON -40.500000  48.460000 -39.660000  48.460000 -39.660000  47.620000 ;
        POLYGON -40.200000  22.685000 -37.845000  20.330000 -40.200000  20.330000 ;
        POLYGON -40.175000 122.495000 -40.175000 120.650000 -42.020000 120.650000 ;
        POLYGON -40.015000  36.655000 -37.665000  36.655000 -37.665000  34.305000 ;
        POLYGON -39.695000 115.980000 -38.210000 115.980000 -39.695000 114.495000 ;
        POLYGON -39.660000  47.620000 -37.660000  47.620000 -37.660000  45.620000 ;
        POLYGON -39.660000 100.370000 -39.660000  99.530000 -40.500000  99.530000 ;
        POLYGON -39.660000 111.690000 -39.660000 108.850000 -42.500000 108.850000 ;
        POLYGON -39.535000 100.495000 -39.535000 100.370000 -39.660000 100.370000 ;
        POLYGON -39.535000 105.530000 -37.340000 105.530000 -39.535000 103.335000 ;
        POLYGON -39.180000  44.300000 -36.375000  41.495000 -39.180000  41.495000 ;
        POLYGON -39.135000  24.455000 -37.365000  24.455000 -37.365000  22.685000 ;
        POLYGON -38.820000 146.495000 -38.820000 138.495000 -46.820000 138.495000 ;
        POLYGON -38.690000 135.295000 -38.690000 132.445000 -41.540000 132.445000 ;
        POLYGON -38.640000  12.645000 -38.340000  12.645000 -38.340000  12.345000 ;
        POLYGON -38.340000   9.495000 -36.340000   7.495000 -38.340000   7.495000 ;
        POLYGON -38.340000  12.345000 -35.490000  12.345000 -35.490000   9.495000 ;
        POLYGON -38.340000 140.495000 -36.340000 140.495000 -38.340000 138.495000 ;
        POLYGON -38.210000 118.815000 -35.375000 118.815000 -38.210000 115.980000 ;
        POLYGON -38.210000 127.660000 -37.845000 127.660000 -38.210000 127.295000 ;
        POLYGON -38.210000 135.775000 -38.210000 135.295000 -38.690000 135.295000 ;
        POLYGON -38.175000 124.495000 -38.175000 122.495000 -40.175000 122.495000 ;
        POLYGON -37.845000  20.330000 -35.010000  17.495000 -37.845000  17.495000 ;
        POLYGON -37.845000 130.495000 -35.010000 130.495000 -37.845000 127.660000 ;
        POLYGON -37.695000  31.495000 -34.855000  28.655000 -37.695000  28.655000 ;
        POLYGON -37.665000  34.305000 -34.855000  34.305000 -34.855000  31.495000 ;
        POLYGON -37.660000  45.620000 -36.340000  45.620000 -36.340000  44.300000 ;
        POLYGON -37.660000 102.370000 -37.660000 100.495000 -39.535000 100.495000 ;
        POLYGON -37.365000  22.685000 -35.010000  22.685000 -35.010000  20.330000 ;
        POLYGON -37.340000 107.535000 -35.335000 107.535000 -37.340000 105.530000 ;
        POLYGON -36.855000 114.495000 -36.855000 111.690000 -39.660000 111.690000 ;
        POLYGON -36.695000 103.335000 -36.695000 102.370000 -37.660000 102.370000 ;
        POLYGON -36.375000  41.495000 -34.375000  39.495000 -36.375000  39.495000 ;
        POLYGON -36.340000  44.300000 -33.535000  44.300000 -33.535000  41.495000 ;
        POLYGON -35.490000 138.495000 -35.490000 135.775000 -38.210000 135.775000 ;
        POLYGON -35.375000 120.650000 -33.540000 120.650000 -35.375000 118.815000 ;
        POLYGON -35.375000 127.295000 -35.375000 124.495000 -38.175000 124.495000 ;
        POLYGON -35.370000 115.980000 -35.370000 114.495000 -36.855000 114.495000 ;
        POLYGON -35.335000 110.335000 -32.535000 110.335000 -35.335000 107.535000 ;
        POLYGON -35.010000  17.495000 -33.010000  15.495000 -35.010000  15.495000 ;
        POLYGON -35.010000  20.330000 -32.175000  20.330000 -32.175000  17.495000 ;
        POLYGON -35.010000 127.660000 -35.010000 127.295000 -35.375000 127.295000 ;
        POLYGON -35.010000 132.495000 -33.010000 132.495000 -35.010000 130.495000 ;
        POLYGON -34.855000  28.655000 -34.535000  28.335000 -34.855000  28.335000 ;
        POLYGON -34.855000  31.495000 -32.015000  31.495000 -32.015000  28.655000 ;
        POLYGON -34.535000  28.335000 -31.695000  25.495000 -34.535000  25.495000 ;
        POLYGON -34.500000  50.940000 -32.500000  48.940000 -34.500000  48.940000 ;
        POLYGON -34.500000  99.050000 -32.500000  99.050000 -34.500000  97.050000 ;
        POLYGON -34.500000 105.530000 -34.500000 103.335000 -36.695000 103.335000 ;
        POLYGON -34.375000  39.495000 -31.535000  36.655000 -34.375000  36.655000 ;
        POLYGON -33.540000 121.685000 -32.505000 121.685000 -33.540000 120.650000 ;
        POLYGON -33.535000  41.495000 -31.535000  41.495000 -31.535000  39.495000 ;
        POLYGON -32.535000 112.170000 -30.700000 112.170000 -32.535000 110.335000 ;
        POLYGON -32.535000 118.815000 -32.535000 115.980000 -35.370000 115.980000 ;
        POLYGON -32.505000 124.495000 -29.695000 124.495000 -32.505000 121.685000 ;
        POLYGON -32.500000  48.940000 -31.055000  47.495000 -32.500000  47.495000 ;
        POLYGON -32.500000  51.780000 -31.660000  51.780000 -31.660000  50.940000 ;
        POLYGON -32.500000 100.495000 -31.055000 100.495000 -32.500000  99.050000 ;
        POLYGON -32.495000 107.535000 -32.495000 105.530000 -34.500000 105.530000 ;
        POLYGON -32.175000 130.495000 -32.175000 127.660000 -35.010000 127.660000 ;
        POLYGON -32.015000  28.655000 -31.695000  28.655000 -31.695000  28.335000 ;
        POLYGON -31.695000  25.495000 -29.695000  23.495000 -31.695000  23.495000 ;
        POLYGON -31.695000  28.335000 -28.855000  28.335000 -28.855000  25.495000 ;
        POLYGON -31.660000  50.940000 -29.660000  50.940000 -29.660000  48.940000 ;
        POLYGON -31.660000  97.050000 -31.660000  96.210000 -32.500000  96.210000 ;
        POLYGON -31.535000  36.655000 -29.185000  34.305000 -31.535000  34.305000 ;
        POLYGON -31.535000  39.495000 -28.695000  39.495000 -28.695000  36.655000 ;
        POLYGON -31.055000  47.495000 -29.340000  45.780000 -31.055000  45.780000 ;
        POLYGON -31.055000 103.335000 -28.215000 103.335000 -31.055000 100.495000 ;
        POLYGON -30.700000 114.495000 -28.375000 114.495000 -30.700000 112.170000 ;
        POLYGON -30.700000 120.650000 -30.700000 118.815000 -32.535000 118.815000 ;
        POLYGON -29.695000 110.335000 -29.695000 107.535000 -32.495000 107.535000 ;
        POLYGON -29.665000 121.685000 -29.665000 120.650000 -30.700000 120.650000 ;
        POLYGON -29.660000  48.940000 -28.215000  48.940000 -28.215000  47.495000 ;
        POLYGON -29.660000  99.050000 -29.660000  97.050000 -31.660000  97.050000 ;
        POLYGON -29.340000  45.780000 -26.500000  42.940000 -29.340000  42.940000 ;
        POLYGON -29.185000  34.305000 -26.375000  31.495000 -29.185000  31.495000 ;
        POLYGON -28.855000 122.495000 -28.855000 121.685000 -29.665000 121.685000 ;
        POLYGON -28.695000  36.655000 -26.345000  36.655000 -26.345000  34.305000 ;
        POLYGON -28.375000 116.495000 -26.375000 116.495000 -28.375000 114.495000 ;
        POLYGON -28.215000  47.495000 -26.500000  47.495000 -26.500000  45.780000 ;
        POLYGON -28.215000 100.495000 -28.215000  99.050000 -29.660000  99.050000 ;
        POLYGON -28.215000 105.685000 -25.865000 105.685000 -28.215000 103.335000 ;
        POLYGON -27.860000 112.170000 -27.860000 110.335000 -29.695000 110.335000 ;
        POLYGON -26.500000  42.940000 -24.015000  40.455000 -26.500000  40.455000 ;
        POLYGON -26.500000  45.780000 -23.660000  45.780000 -23.660000  42.940000 ;
        POLYGON -26.500000  54.260000 -19.735000  47.495000 -26.500000  47.495000 ;
        POLYGON -26.500000 100.495000 -19.735000 100.495000 -26.500000  93.730000 ;
        POLYGON -26.500000 102.210000 -26.500000 100.495000 -28.215000 100.495000 ;
        POLYGON -26.345000  34.305000 -25.535000  34.305000 -25.535000  33.495000 ;
        POLYGON -25.865000 108.495000 -23.055000 108.495000 -25.865000 105.685000 ;
        POLYGON -25.535000 114.495000 -25.535000 112.170000 -27.860000 112.170000 ;
        POLYGON -25.375000 103.335000 -25.375000 102.210000 -26.500000 102.210000 ;
        POLYGON -24.015000  40.455000 -23.055000  39.495000 -24.015000  39.495000 ;
        POLYGON -23.660000  42.940000 -22.215000  42.940000 -22.215000  41.495000 ;
        POLYGON -23.025000 105.685000 -23.025000 103.335000 -25.375000 103.335000 ;
        POLYGON -22.215000 106.495000 -22.215000 105.685000 -23.025000 105.685000 ;
        POLYGON -13.115000   1.495000  -9.275000   1.495000  -9.275000  -2.345000 ;
        POLYGON  -5.240000 108.495000  -3.240000 108.495000  -3.240000 106.495000 ;
        POLYGON  -5.240000 124.495000  -3.240000 124.495000  -3.240000 122.495000 ;
        POLYGON  -5.240000 140.495000  -3.240000 140.495000  -3.240000 138.495000 ;
        POLYGON  -3.240000  17.495000  -3.240000  15.495000  -5.240000  15.495000 ;
        POLYGON  -3.240000  33.495000  -3.240000  31.495000  -5.240000  31.495000 ;
        POLYGON  -3.240000 106.495000   2.760000 106.495000   2.760000 100.495000 ;
        POLYGON  -3.240000 122.495000   2.760000 122.495000   2.760000 116.495000 ;
        POLYGON  -3.240000 138.495000   2.760000 138.495000   2.760000 132.495000 ;
        POLYGON  -2.760000  15.495000   3.240000  15.495000  -2.760000   9.495000 ;
        POLYGON  -2.760000  31.495000   3.240000  31.495000  -2.760000  25.495000 ;
        POLYGON  -2.760000 114.495000   5.240000 106.495000  -2.760000 106.495000 ;
        POLYGON  -2.760000 130.495000   5.240000 122.495000  -2.760000 122.495000 ;
        POLYGON  -2.760000 146.495000   5.240000 138.495000  -2.760000 138.495000 ;
        POLYGON   2.760000  23.495000   2.760000  17.495000  -3.240000  17.495000 ;
        POLYGON   2.760000  39.495000   2.760000  33.495000  -3.240000  33.495000 ;
        POLYGON   3.240000  17.495000   5.240000  17.495000   3.240000  15.495000 ;
        POLYGON   3.240000  33.495000   5.240000  33.495000   3.240000  31.495000 ;
        POLYGON   9.275000   1.495000  13.115000   1.495000   9.275000  -2.345000 ;
        POLYGON  19.735000 100.495000  26.500000 100.495000  26.500000  93.730000 ;
        POLYGON  22.215000  42.460000  23.180000  42.460000  22.215000  41.495000 ;
        POLYGON  22.215000 106.495000  25.020000 103.690000  22.215000 103.690000 ;
        POLYGON  23.055000 108.495000  25.055000 108.495000  25.055000 106.495000 ;
        POLYGON  23.180000  44.655000  25.375000  44.655000  23.180000  42.460000 ;
        POLYGON  23.535000  39.975000  23.535000  39.495000  23.055000  39.495000 ;
        POLYGON  24.015000  40.455000  24.015000  39.975000  23.535000  39.975000 ;
        POLYGON  25.020000 103.690000  26.500000 102.210000  25.020000 102.210000 ;
        POLYGON  25.055000  41.495000  25.055000  40.455000  24.015000  40.455000 ;
        POLYGON  25.055000 106.495000  27.860000 106.495000  27.860000 103.690000 ;
        POLYGON  25.375000  47.495000  28.215000  47.495000  25.375000  44.655000 ;
        POLYGON  25.535000  35.820000  27.860000  35.820000  25.535000  33.495000 ;
        POLYGON  25.535000 114.495000  27.860000 112.170000  25.535000 112.170000 ;
        POLYGON  26.020000  42.460000  26.020000  41.495000  25.055000  41.495000 ;
        POLYGON  26.375000 116.495000  28.375000 116.495000  28.375000 114.495000 ;
        POLYGON  26.500000  54.260000  26.500000  47.495000  19.735000  47.495000 ;
        POLYGON  26.500000 102.210000  28.695000 100.015000  26.500000 100.015000 ;
        POLYGON  27.860000  36.655000  28.695000  36.655000  27.860000  35.820000 ;
        POLYGON  27.860000 103.690000  29.340000 103.690000  29.340000 102.210000 ;
        POLYGON  27.860000 112.170000  29.695000 110.335000  27.860000 110.335000 ;
        POLYGON  28.215000  44.655000  28.215000  42.460000  26.020000  42.460000 ;
        POLYGON  28.215000  48.940000  29.660000  48.940000  28.215000  47.495000 ;
        POLYGON  28.375000  33.495000  28.375000  31.495000  26.375000  31.495000 ;
        POLYGON  28.375000 114.495000  30.700000 114.495000  30.700000 112.170000 ;
        POLYGON  28.695000  39.140000  31.180000  39.140000  28.695000  36.655000 ;
        POLYGON  28.695000 100.015000  29.660000  99.050000  28.695000  99.050000 ;
        POLYGON  28.855000  27.340000  30.700000  27.340000  28.855000  25.495000 ;
        POLYGON  28.855000 122.495000  31.695000 119.655000  28.855000 119.655000 ;
        POLYGON  29.340000 102.210000  31.535000 102.210000  31.535000 100.015000 ;
        POLYGON  29.660000  51.780000  32.500000  51.780000  29.660000  48.940000 ;
        POLYGON  29.660000  99.050000  32.500000  96.210000  29.660000  96.210000 ;
        POLYGON  29.695000 110.335000  32.495000 107.535000  29.695000 107.535000 ;
        POLYGON  29.695000 124.495000  31.695000 124.495000  31.695000 122.495000 ;
        POLYGON  30.700000  28.655000  32.015000  28.655000  30.700000  27.340000 ;
        POLYGON  30.700000  35.820000  30.700000  33.495000  28.375000  33.495000 ;
        POLYGON  30.700000 112.170000  32.535000 112.170000  32.535000 110.335000 ;
        POLYGON  30.705000  24.505000  30.705000  23.495000  29.695000  23.495000 ;
        POLYGON  31.055000  47.495000  31.055000  44.655000  28.215000  44.655000 ;
        POLYGON  31.180000  41.495000  33.535000  41.495000  31.180000  39.140000 ;
        POLYGON  31.535000  36.655000  31.535000  35.820000  30.700000  35.820000 ;
        POLYGON  31.535000 100.015000  32.500000 100.015000  32.500000  99.050000 ;
        POLYGON  31.695000  25.495000  31.695000  24.505000  30.705000  24.505000 ;
        POLYGON  31.695000 119.655000  32.535000 118.815000  31.695000 118.815000 ;
        POLYGON  31.695000 122.495000  34.535000 122.495000  34.535000 119.655000 ;
        POLYGON  32.015000  31.495000  34.855000  31.495000  32.015000  28.655000 ;
        POLYGON  32.175000  20.330000  35.010000  20.330000  32.175000  17.495000 ;
        POLYGON  32.175000 130.495000  35.010000 127.660000  32.175000 127.660000 ;
        POLYGON  32.495000 107.535000  34.500000 105.530000  32.495000 105.530000 ;
        POLYGON  32.500000  48.940000  32.500000  47.495000  31.055000  47.495000 ;
        POLYGON  32.500000  99.050000  34.500000  99.050000  34.500000  97.050000 ;
        POLYGON  32.535000 110.335000  35.335000 110.335000  35.335000 107.535000 ;
        POLYGON  32.535000 118.815000  35.335000 116.015000  32.535000 116.015000 ;
        POLYGON  33.010000 132.495000  35.010000 132.495000  35.010000 130.495000 ;
        POLYGON  33.535000  44.300000  36.340000  44.300000  33.535000  41.495000 ;
        POLYGON  33.540000  27.340000  33.540000  25.495000  31.695000  25.495000 ;
        POLYGON  34.020000  39.140000  34.020000  36.655000  31.535000  36.655000 ;
        POLYGON  34.500000  50.940000  34.500000  48.940000  32.500000  48.940000 ;
        POLYGON  34.500000 105.530000  37.180000 102.850000  34.500000 102.850000 ;
        POLYGON  34.535000 119.655000  35.375000 119.655000  35.375000 118.815000 ;
        POLYGON  34.855000  28.655000  34.855000  27.340000  33.540000  27.340000 ;
        POLYGON  34.855000  32.935000  36.295000  32.935000  34.855000  31.495000 ;
        POLYGON  35.010000  17.495000  35.010000  15.495000  33.010000  15.495000 ;
        POLYGON  35.010000  20.660000  35.340000  20.660000  35.010000  20.330000 ;
        POLYGON  35.010000 127.660000  37.695000 124.975000  35.010000 124.975000 ;
        POLYGON  35.010000 130.495000  37.845000 130.495000  37.845000 127.660000 ;
        POLYGON  35.335000 107.535000  37.340000 107.535000  37.340000 105.530000 ;
        POLYGON  35.335000 116.015000  36.855000 114.495000  35.335000 114.495000 ;
        POLYGON  35.340000  23.495000  38.175000  23.495000  35.340000  20.660000 ;
        POLYGON  35.375000 118.815000  38.175000 118.815000  38.175000 116.015000 ;
        POLYGON  35.490000  12.215000  38.210000  12.215000  35.490000   9.495000 ;
        POLYGON  35.490000 138.495000  38.340000 135.645000  35.490000 135.645000 ;
        POLYGON  36.295000  35.775000  39.135000  35.775000  36.295000  32.935000 ;
        POLYGON  36.340000  45.620000  37.660000  45.620000  36.340000  44.300000 ;
        POLYGON  36.340000 140.495000  38.340000 140.495000  38.340000 138.495000 ;
        POLYGON  36.375000  41.495000  36.375000  39.140000  34.020000  39.140000 ;
        POLYGON  36.855000 114.495000  39.180000 112.170000  36.855000 112.170000 ;
        POLYGON  37.180000 102.850000  40.015000 100.015000  37.180000 100.015000 ;
        POLYGON  37.340000  42.460000  37.340000  41.495000  36.375000  41.495000 ;
        POLYGON  37.340000 105.530000  40.020000 105.530000  40.020000 102.850000 ;
        POLYGON  37.660000  48.460000  40.500000  48.460000  37.660000  45.620000 ;
        POLYGON  37.695000  31.495000  37.695000  28.655000  34.855000  28.655000 ;
        POLYGON  37.695000 124.975000  40.175000 122.495000  37.695000 122.495000 ;
        POLYGON  37.845000  20.330000  37.845000  17.495000  35.010000  17.495000 ;
        POLYGON  37.845000 127.660000  40.530000 127.660000  40.530000 124.975000 ;
        POLYGON  38.175000  20.660000  38.175000  20.330000  37.845000  20.330000 ;
        POLYGON  38.175000  24.505000  39.185000  24.505000  38.175000  23.495000 ;
        POLYGON  38.175000 116.015000  39.695000 116.015000  39.695000 114.495000 ;
        POLYGON  38.210000  12.695000  38.690000  12.695000  38.210000  12.215000 ;
        POLYGON  38.340000   9.495000  38.340000   7.495000  36.340000   7.495000 ;
        POLYGON  38.340000 135.645000  38.640000 135.345000  38.340000 135.345000 ;
        POLYGON  38.340000 138.495000  41.190000 138.495000  41.190000 135.645000 ;
        POLYGON  38.640000 135.345000  41.490000 132.495000  38.640000 132.495000 ;
        POLYGON  38.690000  15.495000  41.490000  15.495000  38.690000  12.695000 ;
        POLYGON  38.820000   7.495000  44.820000   7.495000  38.820000   1.495000 ;
        POLYGON  38.820000 146.495000  44.820000 140.495000  38.820000 140.495000 ;
        POLYGON  39.135000  32.935000  39.135000  31.495000  37.695000  31.495000 ;
        POLYGON  39.135000  37.655000  41.015000  37.655000  39.135000  35.775000 ;
        POLYGON  39.180000  44.300000  39.180000  42.460000  37.340000  42.460000 ;
        POLYGON  39.180000 112.170000  41.015000 110.335000  39.180000 110.335000 ;
        POLYGON  39.185000  27.340000  42.020000  27.340000  39.185000  24.505000 ;
        POLYGON  39.695000 114.495000  42.020000 114.495000  42.020000 112.170000 ;
        POLYGON  40.015000 100.015000  40.500000  99.530000  40.015000  99.530000 ;
        POLYGON  40.020000 102.850000  42.500000 102.850000  42.500000 100.370000 ;
        POLYGON  40.175000 122.495000  41.985000 120.685000  40.175000 120.685000 ;
        POLYGON  40.500000  45.620000  40.500000  44.300000  39.180000  44.300000 ;
        POLYGON  40.530000 124.975000  43.010000 124.975000  43.010000 122.495000 ;
        POLYGON  41.010000  23.495000  41.010000  20.660000  38.175000  20.660000 ;
        POLYGON  41.015000  40.455000  43.815000  40.455000  41.015000  37.655000 ;
        POLYGON  41.015000 110.335000  43.815000 107.535000  41.015000 107.535000 ;
        POLYGON  41.060000  12.215000  41.060000   9.495000  38.340000   9.495000 ;
        POLYGON  41.190000 135.645000  41.490000 135.645000  41.490000 135.345000 ;
        POLYGON  41.490000  15.975000  41.970000  15.975000  41.490000  15.495000 ;
        POLYGON  41.490000 132.495000  43.490000 130.495000  41.490000 130.495000 ;
        POLYGON  41.490000 135.345000  44.340000 135.345000  44.340000 132.495000 ;
        POLYGON  41.540000  12.695000  41.540000  12.215000  41.060000  12.215000 ;
        POLYGON  41.970000  18.825000  44.820000  18.825000  41.970000  15.975000 ;
        POLYGON  41.975000  35.775000  41.975000  32.935000  39.135000  32.935000 ;
        POLYGON  41.985000 120.685000  44.285000 118.385000  41.985000 118.385000 ;
        POLYGON  42.020000  24.505000  42.020000  23.495000  41.010000  23.495000 ;
        POLYGON  42.020000  29.175000  43.855000  29.175000  42.020000  27.340000 ;
        POLYGON  42.020000 112.170000  43.855000 112.170000  43.855000 110.335000 ;
        POLYGON  42.500000  47.620000  42.500000  45.620000  40.500000  45.620000 ;
        POLYGON  43.010000 122.495000  44.820000 122.495000  44.820000 120.685000 ;
        POLYGON  43.490000 130.495000  44.820000 129.165000  43.490000 129.165000 ;
        POLYGON  43.815000  42.300000  45.660000  42.300000  43.815000  40.455000 ;
        POLYGON  43.815000 107.535000  45.660000 105.690000  43.815000 105.690000 ;
        POLYGON  43.855000  31.495000  46.175000  31.495000  43.855000  29.175000 ;
        POLYGON  43.855000  37.655000  43.855000  35.775000  41.975000  35.775000 ;
        POLYGON  43.855000 110.335000  46.655000 110.335000  46.655000 107.535000 ;
        POLYGON  44.285000 118.385000  46.655000 116.015000  44.285000 116.015000 ;
        POLYGON  44.340000  15.495000  44.340000  12.695000  41.540000  12.695000 ;
        POLYGON  44.340000 132.495000  44.820000 132.495000  44.820000 132.015000 ;
        POLYGON  44.820000  12.215000  49.540000  12.215000  44.820000   7.495000 ;
        POLYGON  44.820000  15.975000  44.820000  15.495000  44.340000  15.495000 ;
        POLYGON  44.820000  21.175000  47.170000  21.175000  44.820000  18.825000 ;
        POLYGON  44.820000 120.685000  47.120000 120.685000  47.120000 118.385000 ;
        POLYGON  44.820000 129.165000  47.120000 126.865000  44.820000 126.865000 ;
        POLYGON  44.820000 132.015000  46.340000 132.015000  46.340000 130.495000 ;
        POLYGON  44.820000 140.495000  53.300000 132.015000  44.820000 132.015000 ;
        POLYGON  44.855000  27.340000  44.855000  24.505000  42.020000  24.505000 ;
        POLYGON  45.660000  45.140000  48.500000  45.140000  45.660000  42.300000 ;
        POLYGON  45.660000 105.690000  48.500000 102.850000  45.660000 102.850000 ;
        POLYGON  46.175000  32.985000  47.665000  32.985000  46.175000  31.495000 ;
        POLYGON  46.340000 130.495000  47.670000 130.495000  47.670000 129.165000 ;
        POLYGON  46.655000  40.455000  46.655000  37.655000  43.855000  37.655000 ;
        POLYGON  46.655000 107.535000  48.500000 107.535000  48.500000 105.690000 ;
        POLYGON  46.655000 116.015000  48.175000 114.495000  46.655000 114.495000 ;
        POLYGON  46.690000  29.175000  46.690000  27.340000  44.855000  27.340000 ;
        POLYGON  47.120000 118.385000  49.490000 118.385000  49.490000 116.015000 ;
        POLYGON  47.120000 126.865000  49.970000 124.015000  47.120000 124.015000 ;
        POLYGON  47.170000  24.025000  50.020000  24.025000  47.170000  21.175000 ;
        POLYGON  47.665000  35.775000  50.455000  35.775000  47.665000  32.985000 ;
        POLYGON  47.670000  18.825000  47.670000  15.975000  44.820000  15.975000 ;
        POLYGON  47.670000 129.165000  49.970000 129.165000  49.970000 126.865000 ;
        POLYGON  48.175000 114.495000  50.500000 112.170000  48.175000 112.170000 ;
        POLYGON  48.500000  42.300000  48.500000  40.455000  46.655000  40.455000 ;
        POLYGON  48.500000 105.690000  50.500000 105.690000  50.500000 103.690000 ;
        POLYGON  49.010000  31.495000  49.010000  29.175000  46.690000  29.175000 ;
        POLYGON  49.490000 116.015000  51.010000 116.015000  51.010000 114.495000 ;
        POLYGON  49.540000  18.825000  56.150000  18.825000  49.540000  12.215000 ;
        POLYGON  49.970000 124.015000  51.490000 122.495000  49.970000 122.495000 ;
        POLYGON  49.970000 126.865000  52.820000 126.865000  52.820000 124.015000 ;
        POLYGON  50.020000  21.175000  50.020000  18.825000  47.670000  18.825000 ;
        POLYGON  50.020000  24.455000  50.450000  24.455000  50.020000  24.025000 ;
        POLYGON  50.450000  27.305000  53.300000  27.305000  50.450000  24.455000 ;
        POLYGON  50.450000  32.935000  50.450000  31.495000  49.010000  31.495000 ;
        POLYGON  50.455000  36.655000  51.335000  36.655000  50.455000  35.775000 ;
        POLYGON  50.500000  32.985000  50.500000  32.935000  50.450000  32.935000 ;
        POLYGON  50.500000  44.300000  50.500000  42.300000  48.500000  42.300000 ;
        POLYGON  50.500000 112.170000  53.185000 109.485000  50.500000 109.485000 ;
        POLYGON  51.010000 114.495000  53.335000 114.495000  53.335000 112.170000 ;
        POLYGON  51.335000  38.985000  53.665000  38.985000  51.335000  36.655000 ;
        POLYGON  51.490000 122.495000  53.300000 120.685000  51.490000 120.685000 ;
        POLYGON  52.820000 124.015000  53.300000 124.015000  53.300000 123.535000 ;
        POLYGON  52.870000  24.025000  52.870000  21.175000  50.020000  21.175000 ;
        POLYGON  53.185000 109.485000  55.665000 107.005000  53.185000 107.005000 ;
        POLYGON  53.290000  35.775000  53.290000  32.985000  50.500000  32.985000 ;
        POLYGON  53.300000  24.455000  53.300000  24.025000  52.870000  24.025000 ;
        POLYGON  53.300000  29.655000  55.650000  29.655000  53.300000  27.305000 ;
        POLYGON  53.300000 120.685000  55.600000 118.385000  53.300000 118.385000 ;
        POLYGON  53.300000 123.535000  54.340000 123.535000  54.340000 122.495000 ;
        POLYGON  53.300000 132.015000  61.780000 123.535000  53.300000 123.535000 ;
        POLYGON  53.335000 112.170000  56.020000 112.170000  56.020000 109.485000 ;
        POLYGON  53.665000  41.820000  56.500000  41.820000  53.665000  38.985000 ;
        POLYGON  54.170000  36.655000  54.170000  35.775000  53.290000  35.775000 ;
        POLYGON  54.340000 122.495000  56.150000 122.495000  56.150000 120.685000 ;
        POLYGON  55.600000 118.385000  58.450000 115.535000  55.600000 115.535000 ;
        POLYGON  55.650000  32.505000  58.500000  32.505000  55.650000  29.655000 ;
        POLYGON  55.665000 107.005000  56.500000 106.170000  55.665000 106.170000 ;
        POLYGON  56.020000 109.485000  58.500000 109.485000  58.500000 107.005000 ;
        POLYGON  56.150000  27.305000  56.150000  24.455000  53.300000  24.455000 ;
        POLYGON  56.150000  27.305000  64.630000  27.305000  56.150000  18.825000 ;
        POLYGON  56.150000 120.685000  58.450000 120.685000  58.450000 118.385000 ;
        POLYGON  56.500000  38.985000  56.500000  36.655000  54.170000  36.655000 ;
        POLYGON  58.450000 115.535000  58.980000 115.005000  58.450000 115.005000 ;
        POLYGON  58.450000 118.385000  61.300000 118.385000  61.300000 115.535000 ;
        POLYGON  58.500000  29.655000  58.500000  27.305000  56.150000  27.305000 ;
        POLYGON  58.500000  32.935000  58.930000  32.935000  58.500000  32.505000 ;
        POLYGON  58.500000  40.985000  58.500000  38.985000  56.500000  38.985000 ;
        POLYGON  58.930000  35.655000  61.650000  35.655000  58.930000  32.935000 ;
        POLYGON  58.980000 115.005000  61.770000 112.215000  58.980000 112.215000 ;
        POLYGON  61.300000 115.535000  61.780000 115.535000  61.780000 115.055000 ;
        POLYGON  61.350000  32.505000  61.350000  29.655000  58.500000  29.655000 ;
        POLYGON  61.650000  38.505000  64.500000  38.505000  61.650000  35.655000 ;
        POLYGON  61.770000 112.215000  64.500000 109.485000  61.770000 109.485000 ;
        POLYGON  61.780000  32.935000  61.780000  32.505000  61.350000  32.505000 ;
        POLYGON  61.780000 115.055000  61.830000 115.055000  61.830000 115.005000 ;
        POLYGON  61.780000 123.535000  70.260000 115.055000  61.780000 115.055000 ;
        POLYGON  61.830000 115.005000  64.620000 115.005000  64.620000 112.215000 ;
        POLYGON  64.500000  35.655000  64.500000  32.935000  61.780000  32.935000 ;
        POLYGON  64.620000 112.215000  66.500000 112.215000  66.500000 110.335000 ;
        POLYGON  64.630000  35.175000  72.500000  35.175000  64.630000  27.305000 ;
        POLYGON  66.500000  37.655000  66.500000  35.655000  64.500000  35.655000 ;
        POLYGON  70.260000 115.055000  72.500000 112.815000  70.260000 112.815000 ;
        RECT -72.500000  35.175000 -64.500000  35.655000 ;
        RECT -72.500000  35.655000 -66.500000 112.635000 ;
        RECT -72.500000 112.635000 -64.200000 112.815000 ;
        RECT -69.335000 112.815000 -64.200000 115.485000 ;
        RECT -69.335000 115.485000 -61.350000 115.980000 ;
        RECT -64.615000  27.290000 -57.985000  29.140000 ;
        RECT -64.615000  29.140000 -60.340000  31.495000 ;
        RECT -64.615000  31.495000 -61.780000  32.935000 ;
        RECT -64.615000  32.935000 -64.500000  35.175000 ;
        RECT -64.500000  38.505000 -56.500000  38.985000 ;
        RECT -64.500000  38.985000 -58.500000 107.535000 ;
        RECT -64.500000 107.535000 -57.970000 109.485000 ;
        RECT -63.650000  37.655000 -56.500000  38.505000 ;
        RECT -63.650000 109.485000 -57.970000 110.335000 ;
        RECT -61.650000  35.655000 -55.170000  37.655000 ;
        RECT -61.350000 110.335000 -55.170000 112.170000 ;
        RECT -61.350000 112.170000 -53.335000 112.635000 ;
        RECT -61.350000 118.335000 -58.500000 121.115000 ;
        RECT -61.350000 121.115000 -55.720000 123.965000 ;
        RECT -58.930000  32.935000 -53.170000  35.655000 ;
        RECT -58.500000 112.635000 -53.335000 115.005000 ;
        RECT -58.500000 115.005000 -50.500000 115.485000 ;
        RECT -57.655000  20.330000 -51.530000  22.685000 ;
        RECT -57.655000  22.685000 -53.300000  24.455000 ;
        RECT -57.655000  24.455000 -56.135000  27.290000 ;
        RECT -57.490000  31.495000 -50.450000  32.935000 ;
        RECT -56.500000  41.820000 -48.500000  42.300000 ;
        RECT -56.500000  42.300000 -50.500000 106.170000 ;
        RECT -55.665000  40.985000 -48.500000  41.820000 ;
        RECT -55.665000 106.170000 -48.020000 107.005000 ;
        RECT -55.650000 115.485000 -50.500000 115.980000 ;
        RECT -55.650000 115.980000 -49.525000 118.335000 ;
        RECT -55.135000  29.140000 -49.010000  31.495000 ;
        RECT -55.135000 107.005000 -48.020000 107.535000 ;
        RECT -53.665000  38.985000 -45.695000  39.495000 ;
        RECT -53.665000  39.495000 -48.500000  40.985000 ;
        RECT -53.285000  27.290000 -46.655000  29.140000 ;
        RECT -52.870000 118.335000 -49.525000 118.815000 ;
        RECT -52.870000 118.815000 -46.690000 120.650000 ;
        RECT -52.870000 120.650000 -44.855000 121.115000 ;
        RECT -52.870000 126.815000 -50.020000 129.595000 ;
        RECT -52.870000 129.595000 -47.240000 132.445000 ;
        RECT -52.820000  15.495000 -46.340000  17.495000 ;
        RECT -52.820000  17.495000 -49.175000  20.330000 ;
        RECT -52.335000  37.655000 -45.695000  38.985000 ;
        RECT -52.335000 107.535000 -48.020000 108.850000 ;
        RECT -52.335000 108.850000 -45.340000 110.335000 ;
        RECT -50.500000 110.335000 -45.340000 111.690000 ;
        RECT -50.500000 111.690000 -42.500000 112.170000 ;
        RECT -50.450000  24.455000 -44.805000  27.290000 ;
        RECT -50.335000  35.655000 -42.855000  36.655000 ;
        RECT -50.335000  36.655000 -45.695000  37.655000 ;
        RECT -50.020000 121.115000 -44.855000 122.495000 ;
        RECT -50.020000 122.495000 -43.010000 123.965000 ;
        RECT -49.540000 132.445000 -44.390000 135.295000 ;
        RECT -49.540000 135.295000 -41.540000 135.775000 ;
        RECT -48.680000  22.685000 -41.970000  24.455000 ;
        RECT -48.500000  45.140000 -40.500000  45.620000 ;
        RECT -48.500000  45.620000 -42.500000 100.495000 ;
        RECT -48.500000 100.495000 -42.375000 102.850000 ;
        RECT -48.015000 102.850000 -42.375000 103.335000 ;
        RECT -47.665000 112.170000 -42.500000 114.495000 ;
        RECT -47.665000 114.495000 -39.695000 115.005000 ;
        RECT -47.660000  44.300000 -40.500000  45.140000 ;
        RECT -47.660000 103.335000 -39.535000 103.690000 ;
        RECT -47.615000  32.935000 -40.505000  34.305000 ;
        RECT -47.615000  34.305000 -42.855000  35.655000 ;
        RECT -47.170000 123.965000 -43.010000 124.495000 ;
        RECT -47.170000 124.495000 -41.010000 126.815000 ;
        RECT -46.820000 135.775000 -41.060000 138.495000 ;
        RECT -46.690000 115.005000 -39.695000 115.980000 ;
        RECT -46.325000  20.330000 -40.200000  22.685000 ;
        RECT -46.175000  31.495000 -40.505000  32.935000 ;
        RECT -45.660000  42.300000 -39.180000  44.300000 ;
        RECT -45.180000 103.690000 -39.535000 105.530000 ;
        RECT -45.180000 105.530000 -37.340000 106.170000 ;
        RECT -44.820000   7.495000 -38.340000   9.495000 ;
        RECT -44.820000   9.495000 -41.190000  12.345000 ;
        RECT -44.820000  12.345000 -41.490000  12.645000 ;
        RECT -44.820000  12.645000 -44.340000  15.495000 ;
        RECT -44.390000 126.815000 -41.010000 127.295000 ;
        RECT -44.390000 127.295000 -38.210000 127.660000 ;
        RECT -44.390000 127.660000 -37.845000 129.595000 ;
        RECT -43.855000 115.980000 -38.210000 118.815000 ;
        RECT -43.820000  29.140000 -37.695000  31.495000 ;
        RECT -43.490000  17.495000 -37.845000  20.330000 ;
        RECT -42.855000  39.495000 -36.375000  41.495000 ;
        RECT -42.855000  41.495000 -39.180000  42.300000 ;
        RECT -42.855000 106.170000 -37.340000 107.535000 ;
        RECT -42.855000 107.535000 -35.335000 108.495000 ;
        RECT -42.500000 108.495000 -35.335000 108.850000 ;
        RECT -42.020000 118.815000 -35.375000 120.650000 ;
        RECT -41.970000  27.290000 -34.535000  28.335000 ;
        RECT -41.970000  28.335000 -34.855000  28.655000 ;
        RECT -41.970000  28.655000 -37.695000  29.140000 ;
        RECT -41.540000 129.595000 -37.845000 130.495000 ;
        RECT -41.540000 130.495000 -35.010000 132.445000 ;
        RECT -41.490000  15.495000 -35.010000  17.495000 ;
        RECT -40.500000  48.460000 -32.500000  48.940000 ;
        RECT -40.500000  48.940000 -34.500000  99.050000 ;
        RECT -40.500000  99.050000 -32.500000  99.530000 ;
        RECT -40.175000 120.650000 -33.540000 121.685000 ;
        RECT -40.175000 121.685000 -32.505000 122.495000 ;
        RECT -40.015000  36.655000 -34.375000  39.495000 ;
        RECT -39.660000  47.620000 -32.500000  48.460000 ;
        RECT -39.660000  99.530000 -32.500000 100.370000 ;
        RECT -39.660000 108.850000 -35.335000 110.335000 ;
        RECT -39.660000 110.335000 -32.535000 111.690000 ;
        RECT -39.535000 100.370000 -32.500000 100.495000 ;
        RECT -39.135000  24.455000 -31.695000  25.495000 ;
        RECT -39.135000  25.495000 -34.535000  27.290000 ;
        RECT -38.820000   1.495000  -6.275000   7.495000 ;
        RECT -38.820000 138.495000 -38.340000 140.495000 ;
        RECT -38.820000 140.495000  -2.760000 146.495000 ;
        RECT -38.690000 132.445000 -35.010000 132.495000 ;
        RECT -38.690000 132.495000  -6.080000 135.295000 ;
        RECT -38.640000  12.645000  -2.760000  15.495000 ;
        RECT -38.340000  12.345000  -2.760000  12.645000 ;
        RECT -38.210000 135.295000  -6.080000 135.775000 ;
        RECT -38.175000 122.495000 -32.505000 124.495000 ;
        RECT -37.665000  34.305000 -31.535000  36.655000 ;
        RECT -37.660000  45.620000 -29.340000  45.780000 ;
        RECT -37.660000  45.780000 -31.055000  47.495000 ;
        RECT -37.660000  47.495000 -32.500000  47.620000 ;
        RECT -37.660000 100.495000 -31.055000 102.370000 ;
        RECT -37.365000  22.685000  -6.080000  23.495000 ;
        RECT -37.365000  23.495000 -31.695000  24.455000 ;
        RECT -36.855000 111.690000 -32.535000 112.170000 ;
        RECT -36.855000 112.170000 -30.700000 114.495000 ;
        RECT -36.695000 102.370000 -31.055000 103.335000 ;
        RECT -36.340000  44.300000 -29.340000  45.620000 ;
        RECT -35.490000   9.495000  -2.760000  12.345000 ;
        RECT -35.490000 135.775000  -6.080000 138.495000 ;
        RECT -35.375000 124.495000  -2.760000 127.295000 ;
        RECT -35.370000 114.495000 -28.375000 115.980000 ;
        RECT -35.010000  20.330000  -6.080000  22.685000 ;
        RECT -35.010000 127.295000  -2.760000 127.660000 ;
        RECT -34.855000  31.495000 -29.185000  34.305000 ;
        RECT -34.500000 103.335000 -28.215000 105.530000 ;
        RECT -33.535000  41.495000 -26.500000  42.940000 ;
        RECT -33.535000  42.940000 -29.340000  44.300000 ;
        RECT -32.535000 115.980000 -28.375000 116.495000 ;
        RECT -32.535000 116.495000  -6.080000 118.815000 ;
        RECT -32.500000  51.780000 -26.500000  96.210000 ;
        RECT -32.495000 105.530000 -28.215000 105.685000 ;
        RECT -32.495000 105.685000 -25.865000 107.535000 ;
        RECT -32.175000  17.495000  -6.080000  20.330000 ;
        RECT -32.175000 127.660000  -2.760000 130.495000 ;
        RECT -32.015000  28.655000  -2.760000  31.495000 ;
        RECT -31.695000  28.335000  -2.760000  28.655000 ;
        RECT -31.660000  50.940000 -26.500000  51.780000 ;
        RECT -31.660000  96.210000 -26.500000  97.050000 ;
        RECT -31.535000  39.495000 -24.015000  40.455000 ;
        RECT -31.535000  40.455000 -26.500000  41.495000 ;
        RECT -30.700000 118.815000  -6.080000 120.650000 ;
        RECT -29.695000 107.535000 -25.865000 108.495000 ;
        RECT -29.695000 108.495000  -2.760000 110.335000 ;
        RECT -29.665000 120.650000  -6.080000 121.685000 ;
        RECT -29.660000  48.940000 -26.500000  50.940000 ;
        RECT -29.660000  97.050000 -26.500000  99.050000 ;
        RECT -28.855000  25.495000  -2.760000  28.335000 ;
        RECT -28.855000 121.685000  -6.080000 122.495000 ;
        RECT -28.695000  36.655000  -6.080000  39.495000 ;
        RECT -28.215000  47.495000 -26.500000  48.940000 ;
        RECT -28.215000  99.050000 -26.500000 100.495000 ;
        RECT -27.860000 110.335000  -2.760000 112.170000 ;
        RECT -26.500000  45.780000  25.375000  47.495000 ;
        RECT -26.500000 100.495000  -6.080000 102.210000 ;
        RECT -26.345000  34.305000  -6.080000  36.655000 ;
        RECT -25.535000  33.495000  -6.080000  34.305000 ;
        RECT -25.535000 112.170000  -2.760000 114.495000 ;
        RECT -25.375000 102.210000  -6.080000 103.335000 ;
        RECT -23.660000  42.940000  23.180000  44.655000 ;
        RECT -23.660000  44.655000  25.375000  45.780000 ;
        RECT -23.025000 103.335000  -6.080000 105.685000 ;
        RECT -22.215000  41.495000  22.215000  42.460000 ;
        RECT -22.215000  42.460000  23.180000  42.940000 ;
        RECT -22.215000 105.685000  -6.080000 106.495000 ;
        RECT  -9.275000  -5.950000  -6.275000   1.495000 ;
        RECT  -3.240000  15.495000   3.240000  17.495000 ;
        RECT  -3.240000  31.495000   3.240000  33.495000 ;
        RECT  -3.240000 106.495000  -2.760000 108.495000 ;
        RECT  -3.240000 122.495000  -2.760000 124.495000 ;
        RECT  -3.240000 138.495000  -2.760000 140.495000 ;
        RECT   2.760000  17.495000  32.175000  20.330000 ;
        RECT   2.760000  20.330000  35.010000  20.660000 ;
        RECT   2.760000  20.660000  35.340000  23.495000 ;
        RECT   2.760000  33.495000  25.535000  35.820000 ;
        RECT   2.760000  35.820000  27.860000  36.655000 ;
        RECT   2.760000  36.655000  28.695000  39.140000 ;
        RECT   2.760000  39.140000  31.180000  39.495000 ;
        RECT   2.760000 100.495000  26.500000 102.210000 ;
        RECT   2.760000 102.210000  25.020000 103.690000 ;
        RECT   2.760000 103.690000  22.215000 106.495000 ;
        RECT   2.760000 116.495000  32.535000 118.815000 ;
        RECT   2.760000 118.815000  31.695000 119.655000 ;
        RECT   2.760000 119.655000  28.855000 122.495000 ;
        RECT   2.760000 132.495000  38.640000 135.345000 ;
        RECT   2.760000 135.345000  38.340000 135.645000 ;
        RECT   2.760000 135.645000  35.490000 138.495000 ;
        RECT   6.080000   9.495000  35.490000  12.215000 ;
        RECT   6.080000  12.215000  38.210000  12.695000 ;
        RECT   6.080000  12.695000  38.690000  15.495000 ;
        RECT   6.080000  25.495000  28.855000  27.340000 ;
        RECT   6.080000  27.340000  30.700000  28.655000 ;
        RECT   6.080000  28.655000  32.015000  31.495000 ;
        RECT   6.080000 108.495000  29.695000 110.335000 ;
        RECT   6.080000 110.335000  27.860000 112.170000 ;
        RECT   6.080000 112.170000  25.535000 114.495000 ;
        RECT   6.080000 124.495000  37.695000 124.975000 ;
        RECT   6.080000 124.975000  35.010000 127.660000 ;
        RECT   6.080000 127.660000  32.175000 130.495000 ;
        RECT   6.080000 140.495000  38.820000 146.495000 ;
        RECT   6.275000  -5.950000   9.275000   1.495000 ;
        RECT   6.275000   1.495000  38.820000   7.495000 ;
        RECT  23.535000  39.495000  31.180000  39.975000 ;
        RECT  24.015000  39.975000  31.180000  40.455000 ;
        RECT  25.055000  40.455000  31.180000  41.495000 ;
        RECT  25.055000 106.495000  32.495000 107.535000 ;
        RECT  25.055000 107.535000  29.695000 108.495000 ;
        RECT  26.020000  41.495000  33.535000  42.460000 ;
        RECT  26.500000  47.495000  28.215000  48.940000 ;
        RECT  26.500000  48.940000  29.660000  51.780000 ;
        RECT  26.500000  51.780000  32.500000  96.210000 ;
        RECT  26.500000  96.210000  29.660000  99.050000 ;
        RECT  26.500000  99.050000  28.695000 100.015000 ;
        RECT  27.860000 103.690000  34.500000 105.530000 ;
        RECT  27.860000 105.530000  32.495000 106.495000 ;
        RECT  28.215000  42.460000  33.535000  44.300000 ;
        RECT  28.215000  44.300000  36.340000  44.655000 ;
        RECT  28.375000  31.495000  34.855000  32.935000 ;
        RECT  28.375000  32.935000  36.295000  33.495000 ;
        RECT  28.375000 114.495000  35.335000 116.015000 ;
        RECT  28.375000 116.015000  32.535000 116.495000 ;
        RECT  29.340000 102.210000  37.180000 102.850000 ;
        RECT  29.340000 102.850000  34.500000 103.690000 ;
        RECT  30.700000  33.495000  36.295000  35.775000 ;
        RECT  30.700000  35.775000  39.135000  35.820000 ;
        RECT  30.700000 112.170000  36.855000 114.495000 ;
        RECT  30.705000  23.495000  38.175000  24.505000 ;
        RECT  31.055000  44.655000  36.340000  45.620000 ;
        RECT  31.055000  45.620000  37.660000  47.495000 ;
        RECT  31.535000  35.820000  39.135000  36.655000 ;
        RECT  31.535000 100.015000  37.180000 102.210000 ;
        RECT  31.695000  24.505000  39.185000  25.495000 ;
        RECT  31.695000 122.495000  37.695000 124.495000 ;
        RECT  32.500000  47.495000  37.660000  48.460000 ;
        RECT  32.500000  48.460000  40.500000  48.940000 ;
        RECT  32.500000  99.050000  40.500000  99.530000 ;
        RECT  32.500000  99.530000  40.015000 100.015000 ;
        RECT  32.535000 110.335000  39.180000 112.170000 ;
        RECT  33.540000  25.495000  39.185000  27.340000 ;
        RECT  34.020000  36.655000  39.135000  37.655000 ;
        RECT  34.020000  37.655000  41.015000  39.140000 ;
        RECT  34.500000  48.940000  40.500000  99.050000 ;
        RECT  34.535000 119.655000  41.985000 120.685000 ;
        RECT  34.535000 120.685000  40.175000 122.495000 ;
        RECT  34.855000  27.340000  42.020000  28.655000 ;
        RECT  35.010000  15.495000  41.490000  15.975000 ;
        RECT  35.010000  15.975000  41.970000  17.495000 ;
        RECT  35.010000 130.495000  41.490000 132.495000 ;
        RECT  35.335000 107.535000  41.015000 110.335000 ;
        RECT  35.375000 118.815000  41.985000 119.655000 ;
        RECT  36.375000  39.140000  41.015000  40.455000 ;
        RECT  36.375000  40.455000  43.815000  41.495000 ;
        RECT  37.340000  41.495000  43.815000  42.300000 ;
        RECT  37.340000  42.300000  45.660000  42.460000 ;
        RECT  37.340000 105.530000  45.660000 105.690000 ;
        RECT  37.340000 105.690000  43.815000 107.535000 ;
        RECT  37.695000  28.655000  42.020000  29.175000 ;
        RECT  37.695000  29.175000  43.855000  31.495000 ;
        RECT  37.845000  17.495000  41.970000  18.825000 ;
        RECT  37.845000  18.825000  44.820000  20.330000 ;
        RECT  37.845000 127.660000  44.820000 129.165000 ;
        RECT  37.845000 129.165000  43.490000 130.495000 ;
        RECT  38.175000  20.330000  44.820000  20.660000 ;
        RECT  38.175000 116.015000  44.285000 118.385000 ;
        RECT  38.175000 118.385000  41.985000 118.815000 ;
        RECT  38.340000   7.495000  44.820000   9.495000 ;
        RECT  38.340000 138.495000  44.820000 140.495000 ;
        RECT  39.135000  31.495000  46.175000  32.935000 ;
        RECT  39.180000  42.460000  45.660000  44.300000 ;
        RECT  39.695000 114.495000  46.655000 116.015000 ;
        RECT  40.020000 102.850000  45.660000 105.530000 ;
        RECT  40.500000  44.300000  45.660000  45.140000 ;
        RECT  40.500000  45.140000  48.500000  45.620000 ;
        RECT  40.530000 124.975000  47.120000 126.865000 ;
        RECT  40.530000 126.865000  44.820000 127.660000 ;
        RECT  41.010000  20.660000  44.820000  21.175000 ;
        RECT  41.010000  21.175000  47.170000  23.495000 ;
        RECT  41.060000   9.495000  44.820000  12.215000 ;
        RECT  41.190000 135.645000  44.820000 138.495000 ;
        RECT  41.490000 135.345000  44.820000 135.645000 ;
        RECT  41.540000  12.215000  49.540000  12.695000 ;
        RECT  41.975000  32.935000  46.175000  32.985000 ;
        RECT  41.975000  32.985000  47.665000  35.775000 ;
        RECT  42.020000  23.495000  47.170000  24.025000 ;
        RECT  42.020000  24.025000  50.020000  24.455000 ;
        RECT  42.020000  24.455000  50.450000  24.505000 ;
        RECT  42.020000 112.170000  48.175000 114.495000 ;
        RECT  42.500000  45.620000  48.500000 102.850000 ;
        RECT  43.010000 122.495000  49.970000 124.015000 ;
        RECT  43.010000 124.015000  47.120000 124.975000 ;
        RECT  43.855000  35.775000  50.455000  36.655000 ;
        RECT  43.855000  36.655000  51.335000  37.655000 ;
        RECT  43.855000 110.335000  50.500000 112.170000 ;
        RECT  44.340000  12.695000  49.540000  15.495000 ;
        RECT  44.340000 132.495000  44.820000 135.345000 ;
        RECT  44.820000  15.495000  49.540000  15.975000 ;
        RECT  44.820000 120.685000  51.490000 122.495000 ;
        RECT  44.855000  24.505000  50.450000  27.305000 ;
        RECT  44.855000  27.305000  53.300000  27.340000 ;
        RECT  46.340000 130.495000  53.300000 132.015000 ;
        RECT  46.655000  37.655000  51.335000  38.985000 ;
        RECT  46.655000  38.985000  53.665000  40.455000 ;
        RECT  46.655000 107.535000  53.185000 109.485000 ;
        RECT  46.655000 109.485000  50.500000 110.335000 ;
        RECT  46.690000  27.340000  53.300000  29.175000 ;
        RECT  47.120000 118.385000  53.300000 120.685000 ;
        RECT  47.670000  15.975000  49.540000  18.825000 ;
        RECT  47.670000 129.165000  53.300000 130.495000 ;
        RECT  48.500000  40.455000  53.665000  41.820000 ;
        RECT  48.500000  41.820000  56.500000  42.300000 ;
        RECT  48.500000 105.690000  56.500000 106.170000 ;
        RECT  48.500000 106.170000  55.665000 107.005000 ;
        RECT  48.500000 107.005000  53.185000 107.535000 ;
        RECT  49.010000  29.175000  53.300000  29.655000 ;
        RECT  49.010000  29.655000  55.650000  31.495000 ;
        RECT  49.490000 116.015000  55.600000 118.385000 ;
        RECT  49.970000 126.865000  53.300000 129.165000 ;
        RECT  50.020000  18.825000  56.150000  21.175000 ;
        RECT  50.450000  31.495000  55.650000  32.505000 ;
        RECT  50.450000  32.505000  58.500000  32.935000 ;
        RECT  50.500000  32.935000  58.930000  32.985000 ;
        RECT  50.500000  42.300000  56.500000 105.690000 ;
        RECT  51.010000 114.495000  58.980000 115.005000 ;
        RECT  51.010000 115.005000  58.450000 115.535000 ;
        RECT  51.010000 115.535000  55.600000 116.015000 ;
        RECT  52.820000 124.015000  53.300000 126.865000 ;
        RECT  52.870000  21.175000  56.150000  24.025000 ;
        RECT  53.290000  32.985000  58.930000  35.655000 ;
        RECT  53.290000  35.655000  61.650000  35.775000 ;
        RECT  53.300000  24.025000  56.150000  24.455000 ;
        RECT  53.335000 112.170000  61.770000 112.215000 ;
        RECT  53.335000 112.215000  58.980000 114.495000 ;
        RECT  54.170000  35.775000  61.650000  36.655000 ;
        RECT  54.340000 122.495000  61.780000 123.535000 ;
        RECT  56.020000 109.485000  61.770000 112.170000 ;
        RECT  56.150000 120.685000  61.780000 122.495000 ;
        RECT  56.500000  36.655000  61.650000  38.505000 ;
        RECT  56.500000  38.505000  64.500000  38.985000 ;
        RECT  58.450000 118.385000  61.780000 120.685000 ;
        RECT  58.500000  27.305000  64.630000  29.655000 ;
        RECT  58.500000  38.985000  64.500000 109.485000 ;
        RECT  61.300000 115.535000  61.780000 118.385000 ;
        RECT  61.350000  29.655000  64.630000  32.505000 ;
        RECT  61.780000  32.505000  64.630000  32.935000 ;
        RECT  61.830000 115.005000  70.260000 115.055000 ;
        RECT  64.500000  32.935000  64.630000  35.175000 ;
        RECT  64.500000  35.175000  72.500000  35.655000 ;
        RECT  64.620000 112.215000  72.500000 112.815000 ;
        RECT  64.620000 112.815000  70.260000 115.005000 ;
        RECT  66.500000  35.655000  72.500000 112.215000 ;
    END
  END CENTERTAP
  OBS
    LAYER li1 ;
      RECT -98.300000  -8.210000  98.300000  -7.910000 ;
      RECT -98.300000  -7.910000 -98.000000 156.350000 ;
      RECT -98.300000 156.350000  98.300000 156.650000 ;
      RECT -97.000000  -6.630000  97.000000  -5.970000 ;
      RECT -97.000000  -5.410000  97.000000  -4.750000 ;
      RECT -97.000000  -4.190000  97.000000  -3.530000 ;
      RECT -97.000000  -2.970000  97.000000  -2.310000 ;
      RECT -97.000000  -1.750000  97.000000  -1.090000 ;
      RECT -97.000000  -0.530000  97.000000   0.130000 ;
      RECT -97.000000   0.690000  97.000000   1.350000 ;
      RECT -97.000000   1.910000  97.000000   2.570000 ;
      RECT -97.000000   3.130000  97.000000   3.790000 ;
      RECT -97.000000   4.350000  97.000000   5.010000 ;
      RECT -97.000000   5.570000  97.000000   6.230000 ;
      RECT -97.000000   6.790000  97.000000   7.450000 ;
      RECT -97.000000   8.010000  97.000000   8.670000 ;
      RECT -97.000000   9.230000  97.000000   9.890000 ;
      RECT -97.000000  10.450000  97.000000  11.110000 ;
      RECT -97.000000  11.670000  97.000000  12.330000 ;
      RECT -97.000000  12.890000  97.000000  13.550000 ;
      RECT -97.000000  14.110000  97.000000  14.770000 ;
      RECT -97.000000  15.330000  97.000000  15.990000 ;
      RECT -97.000000  16.550000  97.000000  17.210000 ;
      RECT -97.000000  17.770000  97.000000  18.430000 ;
      RECT -97.000000  18.990000  97.000000  19.650000 ;
      RECT -97.000000  20.210000  97.000000  20.870000 ;
      RECT -97.000000  21.430000  97.000000  22.090000 ;
      RECT -97.000000  22.650000  97.000000  23.310000 ;
      RECT -97.000000  23.870000  97.000000  24.530000 ;
      RECT -97.000000  25.090000  97.000000  25.750000 ;
      RECT -97.000000  26.310000  97.000000  26.970000 ;
      RECT -97.000000  27.530000  97.000000  28.190000 ;
      RECT -97.000000  28.750000  97.000000  29.410000 ;
      RECT -97.000000  29.970000  97.000000  30.630000 ;
      RECT -97.000000  31.190000  97.000000  31.850000 ;
      RECT -97.000000  32.410000  97.000000  33.070000 ;
      RECT -97.000000  33.630000  97.000000  34.290000 ;
      RECT -97.000000  34.850000  97.000000  35.510000 ;
      RECT -97.000000  36.070000  97.000000  36.730000 ;
      RECT -97.000000  37.290000  97.000000  37.950000 ;
      RECT -97.000000  38.510000  97.000000  39.170000 ;
      RECT -97.000000  39.730000  97.000000  40.390000 ;
      RECT -97.000000  40.950000  97.000000  41.610000 ;
      RECT -97.000000  42.170000  97.000000  42.830000 ;
      RECT -97.000000  43.390000  97.000000  44.050000 ;
      RECT -97.000000  44.610000  97.000000  45.270000 ;
      RECT -97.000000  45.830000  97.000000  46.490000 ;
      RECT -97.000000  47.050000  97.000000  47.710000 ;
      RECT -97.000000  48.270000  97.000000  48.930000 ;
      RECT -97.000000  49.490000  97.000000  50.150000 ;
      RECT -97.000000  50.710000  97.000000  51.370000 ;
      RECT -97.000000  51.930000  97.000000  52.590000 ;
      RECT -97.000000  53.150000  97.000000  53.810000 ;
      RECT -97.000000  54.370000  97.000000  55.030000 ;
      RECT -97.000000  55.590000  97.000000  56.250000 ;
      RECT -97.000000  56.810000  97.000000  57.470000 ;
      RECT -97.000000  58.030000  97.000000  58.690000 ;
      RECT -97.000000  59.250000  97.000000  59.910000 ;
      RECT -97.000000  60.470000  97.000000  61.130000 ;
      RECT -97.000000  61.690000  97.000000  62.350000 ;
      RECT -97.000000  62.910000  97.000000  63.570000 ;
      RECT -97.000000  64.130000  97.000000  64.790000 ;
      RECT -97.000000  65.350000  97.000000  66.010000 ;
      RECT -97.000000  66.570000  97.000000  67.230000 ;
      RECT -97.000000  67.790000  97.000000  68.450000 ;
      RECT -97.000000  69.010000  97.000000  69.670000 ;
      RECT -97.000000  70.230000  97.000000  70.890000 ;
      RECT -97.000000  71.450000  97.000000  72.110000 ;
      RECT -97.000000  72.670000  97.000000  73.330000 ;
      RECT -97.000000  73.890000  97.000000  74.550000 ;
      RECT -97.000000  75.110000  97.000000  75.770000 ;
      RECT -97.000000  76.330000  97.000000  76.990000 ;
      RECT -97.000000  77.550000  97.000000  78.210000 ;
      RECT -97.000000  78.770000  97.000000  79.430000 ;
      RECT -97.000000  79.990000  97.000000  80.650000 ;
      RECT -97.000000  81.210000  97.000000  81.870000 ;
      RECT -97.000000  82.430000  97.000000  83.090000 ;
      RECT -97.000000  83.650000  97.000000  84.310000 ;
      RECT -97.000000  84.870000  97.000000  85.530000 ;
      RECT -97.000000  86.090000  97.000000  86.750000 ;
      RECT -97.000000  87.310000  97.000000  87.970000 ;
      RECT -97.000000  88.530000  97.000000  89.190000 ;
      RECT -97.000000  89.750000  97.000000  90.410000 ;
      RECT -97.000000  90.970000  97.000000  91.630000 ;
      RECT -97.000000  92.190000  97.000000  92.850000 ;
      RECT -97.000000  93.410000  97.000000  94.070000 ;
      RECT -97.000000  94.630000  97.000000  95.290000 ;
      RECT -97.000000  95.850000  97.000000  96.510000 ;
      RECT -97.000000  97.070000  97.000000  97.730000 ;
      RECT -97.000000  98.290000  97.000000  98.950000 ;
      RECT -97.000000  99.510000  97.000000 100.170000 ;
      RECT -97.000000 100.730000  97.000000 101.390000 ;
      RECT -97.000000 101.950000  97.000000 102.610000 ;
      RECT -97.000000 103.170000  97.000000 103.830000 ;
      RECT -97.000000 104.390000  97.000000 105.050000 ;
      RECT -97.000000 105.610000  97.000000 106.270000 ;
      RECT -97.000000 106.830000  97.000000 107.490000 ;
      RECT -97.000000 108.050000  97.000000 108.710000 ;
      RECT -97.000000 109.270000  97.000000 109.930000 ;
      RECT -97.000000 110.490000  97.000000 111.150000 ;
      RECT -97.000000 111.710000  97.000000 112.370000 ;
      RECT -97.000000 112.930000  97.000000 113.590000 ;
      RECT -97.000000 114.150000  97.000000 114.810000 ;
      RECT -97.000000 115.370000  97.000000 116.030000 ;
      RECT -97.000000 116.590000  97.000000 117.250000 ;
      RECT -97.000000 117.810000  97.000000 118.470000 ;
      RECT -97.000000 119.030000  97.000000 119.690000 ;
      RECT -97.000000 120.250000  97.000000 120.910000 ;
      RECT -97.000000 121.470000  97.000000 122.130000 ;
      RECT -97.000000 122.690000  97.000000 123.350000 ;
      RECT -97.000000 123.910000  97.000000 124.570000 ;
      RECT -97.000000 125.130000  97.000000 125.790000 ;
      RECT -97.000000 126.350000  97.000000 127.010000 ;
      RECT -97.000000 127.570000  97.000000 128.230000 ;
      RECT -97.000000 128.790000  97.000000 129.450000 ;
      RECT -97.000000 130.010000  97.000000 130.670000 ;
      RECT -97.000000 131.230000  97.000000 131.890000 ;
      RECT -97.000000 132.450000  97.000000 133.110000 ;
      RECT -97.000000 133.670000  97.000000 134.330000 ;
      RECT -97.000000 134.890000  97.000000 135.550000 ;
      RECT -97.000000 136.110000  97.000000 136.770000 ;
      RECT -97.000000 137.330000  97.000000 137.990000 ;
      RECT -97.000000 138.550000  97.000000 139.210000 ;
      RECT -97.000000 139.770000  97.000000 140.430000 ;
      RECT -97.000000 140.990000  97.000000 141.650000 ;
      RECT -97.000000 142.210000  97.000000 142.870000 ;
      RECT -97.000000 143.430000  97.000000 144.090000 ;
      RECT -97.000000 144.650000  97.000000 145.310000 ;
      RECT -97.000000 145.870000  97.000000 146.530000 ;
      RECT -97.000000 147.090000  97.000000 147.750000 ;
      RECT -97.000000 148.310000  97.000000 148.970000 ;
      RECT -97.000000 149.530000  97.000000 150.190000 ;
      RECT -97.000000 150.750000  97.000000 151.410000 ;
      RECT -97.000000 151.970000  97.000000 152.630000 ;
      RECT -97.000000 153.190000  97.000000 153.850000 ;
      RECT -97.000000 154.410000  97.000000 155.070000 ;
      RECT  -2.500000  -6.910000   2.500000  -6.630000 ;
      RECT  -2.500000  -5.970000   2.500000  -5.410000 ;
      RECT  -2.500000  -4.750000   2.500000  -4.190000 ;
      RECT  -2.500000  -3.530000   2.500000  -2.970000 ;
      RECT  -2.500000  -2.310000   2.500000  -1.750000 ;
      RECT  -2.500000  -1.090000   2.500000  -0.530000 ;
      RECT  -2.500000   0.130000   2.500000   0.690000 ;
      RECT  -2.500000   1.350000   2.500000   1.910000 ;
      RECT  -2.500000   2.570000   2.500000   3.130000 ;
      RECT  -2.500000   3.790000   2.500000   4.350000 ;
      RECT  -2.500000   5.010000   2.500000   5.570000 ;
      RECT  -2.500000   6.230000   2.500000   6.790000 ;
      RECT  -2.500000   7.450000   2.500000   8.010000 ;
      RECT  -2.500000   8.670000   2.500000   9.230000 ;
      RECT  -2.500000   9.890000   2.500000  10.450000 ;
      RECT  -2.500000  11.110000   2.500000  11.670000 ;
      RECT  -2.500000  12.330000   2.500000  12.890000 ;
      RECT  -2.500000  13.550000   2.500000  14.110000 ;
      RECT  -2.500000  14.770000   2.500000  15.330000 ;
      RECT  -2.500000  15.990000   2.500000  16.550000 ;
      RECT  -2.500000  17.210000   2.500000  17.770000 ;
      RECT  -2.500000  18.430000   2.500000  18.990000 ;
      RECT  -2.500000  19.650000   2.500000  20.210000 ;
      RECT  -2.500000  20.870000   2.500000  21.430000 ;
      RECT  -2.500000  22.090000   2.500000  22.650000 ;
      RECT  -2.500000  23.310000   2.500000  23.870000 ;
      RECT  -2.500000  24.530000   2.500000  25.090000 ;
      RECT  -2.500000  25.750000   2.500000  26.310000 ;
      RECT  -2.500000  26.970000   2.500000  27.530000 ;
      RECT  -2.500000  28.190000   2.500000  28.750000 ;
      RECT  -2.500000  29.410000   2.500000  29.970000 ;
      RECT  -2.500000  30.630000   2.500000  31.190000 ;
      RECT  -2.500000  31.850000   2.500000  32.410000 ;
      RECT  -2.500000  33.070000   2.500000  33.630000 ;
      RECT  -2.500000  34.290000   2.500000  34.850000 ;
      RECT  -2.500000  35.510000   2.500000  36.070000 ;
      RECT  -2.500000  36.730000   2.500000  37.290000 ;
      RECT  -2.500000  37.950000   2.500000  38.510000 ;
      RECT  -2.500000  39.170000   2.500000  39.730000 ;
      RECT  -2.500000  40.390000   2.500000  40.950000 ;
      RECT  -2.500000  41.610000   2.500000  42.170000 ;
      RECT  -2.500000  42.830000   2.500000  43.390000 ;
      RECT  -2.500000  44.050000   2.500000  44.610000 ;
      RECT  -2.500000  45.270000   2.500000  45.830000 ;
      RECT  -2.500000  46.490000   2.500000  47.050000 ;
      RECT  -2.500000  47.710000   2.500000  48.270000 ;
      RECT  -2.500000  48.930000   2.500000  49.490000 ;
      RECT  -2.500000  50.150000   2.500000  50.710000 ;
      RECT  -2.500000  51.370000   2.500000  51.930000 ;
      RECT  -2.500000  52.590000   2.500000  53.150000 ;
      RECT  -2.500000  53.810000   2.500000  54.370000 ;
      RECT  -2.500000  55.030000   2.500000  55.590000 ;
      RECT  -2.500000  56.250000   2.500000  56.810000 ;
      RECT  -2.500000  57.470000   2.500000  58.030000 ;
      RECT  -2.500000  58.690000   2.500000  59.250000 ;
      RECT  -2.500000  59.910000   2.500000  60.470000 ;
      RECT  -2.500000  61.130000   2.500000  61.690000 ;
      RECT  -2.500000  62.350000   2.500000  62.910000 ;
      RECT  -2.500000  63.570000   2.500000  64.130000 ;
      RECT  -2.500000  64.790000   2.500000  65.350000 ;
      RECT  -2.500000  66.010000   2.500000  66.570000 ;
      RECT  -2.500000  67.230000   2.500000  67.790000 ;
      RECT  -2.500000  68.450000   2.500000  69.010000 ;
      RECT  -2.500000  69.670000   2.500000  70.230000 ;
      RECT  -2.500000  70.890000   2.500000  71.450000 ;
      RECT  -2.500000  72.110000   2.500000  72.670000 ;
      RECT  -2.500000  73.330000   2.500000  73.890000 ;
      RECT  -2.500000  74.550000   2.500000  75.110000 ;
      RECT  -2.500000  75.770000   2.500000  76.330000 ;
      RECT  -2.500000  76.990000   2.500000  77.550000 ;
      RECT  -2.500000  78.210000   2.500000  78.770000 ;
      RECT  -2.500000  79.430000   2.500000  79.990000 ;
      RECT  -2.500000  80.650000   2.500000  81.210000 ;
      RECT  -2.500000  81.870000   2.500000  82.430000 ;
      RECT  -2.500000  83.090000   2.500000  83.650000 ;
      RECT  -2.500000  84.310000   2.500000  84.870000 ;
      RECT  -2.500000  85.530000   2.500000  86.090000 ;
      RECT  -2.500000  86.750000   2.500000  87.310000 ;
      RECT  -2.500000  87.970000   2.500000  88.530000 ;
      RECT  -2.500000  89.190000   2.500000  89.750000 ;
      RECT  -2.500000  90.410000   2.500000  90.970000 ;
      RECT  -2.500000  91.630000   2.500000  92.190000 ;
      RECT  -2.500000  92.850000   2.500000  93.410000 ;
      RECT  -2.500000  94.070000   2.500000  94.630000 ;
      RECT  -2.500000  95.290000   2.500000  95.850000 ;
      RECT  -2.500000  96.510000   2.500000  97.070000 ;
      RECT  -2.500000  97.730000   2.500000  98.290000 ;
      RECT  -2.500000  98.950000   2.500000  99.510000 ;
      RECT  -2.500000 100.170000   2.500000 100.730000 ;
      RECT  -2.500000 101.390000   2.500000 101.950000 ;
      RECT  -2.500000 102.610000   2.500000 103.170000 ;
      RECT  -2.500000 103.830000   2.500000 104.390000 ;
      RECT  -2.500000 105.050000   2.500000 105.610000 ;
      RECT  -2.500000 106.270000   2.500000 106.830000 ;
      RECT  -2.500000 107.490000   2.500000 108.050000 ;
      RECT  -2.500000 108.710000   2.500000 109.270000 ;
      RECT  -2.500000 109.930000   2.500000 110.490000 ;
      RECT  -2.500000 111.150000   2.500000 111.710000 ;
      RECT  -2.500000 112.370000   2.500000 112.930000 ;
      RECT  -2.500000 113.590000   2.500000 114.150000 ;
      RECT  -2.500000 114.810000   2.500000 115.370000 ;
      RECT  -2.500000 116.030000   2.500000 116.590000 ;
      RECT  -2.500000 117.250000   2.500000 117.810000 ;
      RECT  -2.500000 118.470000   2.500000 119.030000 ;
      RECT  -2.500000 119.690000   2.500000 120.250000 ;
      RECT  -2.500000 120.910000   2.500000 121.470000 ;
      RECT  -2.500000 122.130000   2.500000 122.690000 ;
      RECT  -2.500000 123.350000   2.500000 123.910000 ;
      RECT  -2.500000 124.570000   2.500000 125.130000 ;
      RECT  -2.500000 125.790000   2.500000 126.350000 ;
      RECT  -2.500000 127.010000   2.500000 127.570000 ;
      RECT  -2.500000 128.230000   2.500000 128.790000 ;
      RECT  -2.500000 129.450000   2.500000 130.010000 ;
      RECT  -2.500000 130.670000   2.500000 131.230000 ;
      RECT  -2.500000 131.890000   2.500000 132.450000 ;
      RECT  -2.500000 133.110000   2.500000 133.670000 ;
      RECT  -2.500000 134.330000   2.500000 134.890000 ;
      RECT  -2.500000 135.550000   2.500000 136.110000 ;
      RECT  -2.500000 136.770000   2.500000 137.330000 ;
      RECT  -2.500000 137.990000   2.500000 138.550000 ;
      RECT  -2.500000 139.210000   2.500000 139.770000 ;
      RECT  -2.500000 140.430000   2.500000 140.990000 ;
      RECT  -2.500000 141.650000   2.500000 142.210000 ;
      RECT  -2.500000 142.870000   2.500000 143.430000 ;
      RECT  -2.500000 144.090000   2.500000 144.650000 ;
      RECT  -2.500000 145.310000   2.500000 145.870000 ;
      RECT  -2.500000 146.530000   2.500000 147.090000 ;
      RECT  -2.500000 147.750000   2.500000 148.310000 ;
      RECT  -2.500000 148.970000   2.500000 149.530000 ;
      RECT  -2.500000 150.190000   2.500000 150.750000 ;
      RECT  -2.500000 151.410000   2.500000 151.970000 ;
      RECT  -2.500000 152.630000   2.500000 153.190000 ;
      RECT  -2.500000 153.850000   2.500000 154.410000 ;
      RECT  -2.500000 155.070000   2.500000 155.350000 ;
      RECT  98.000000  -7.910000  98.300000 156.350000 ;
    LAYER mcon ;
      RECT -98.235000  -7.700000 -98.065000  -7.530000 ;
      RECT -98.235000  -7.340000 -98.065000  -7.170000 ;
      RECT -98.235000  -6.980000 -98.065000  -6.810000 ;
      RECT -98.235000  -6.620000 -98.065000  -6.450000 ;
      RECT -98.235000  -6.260000 -98.065000  -6.090000 ;
      RECT -98.235000  -5.900000 -98.065000  -5.730000 ;
      RECT -98.235000  -5.540000 -98.065000  -5.370000 ;
      RECT -98.235000  -5.180000 -98.065000  -5.010000 ;
      RECT -98.235000  -4.820000 -98.065000  -4.650000 ;
      RECT -98.235000  -4.460000 -98.065000  -4.290000 ;
      RECT -98.235000  -4.100000 -98.065000  -3.930000 ;
      RECT -98.235000  -3.740000 -98.065000  -3.570000 ;
      RECT -98.235000  -3.380000 -98.065000  -3.210000 ;
      RECT -98.235000  -3.020000 -98.065000  -2.850000 ;
      RECT -98.235000  -2.660000 -98.065000  -2.490000 ;
      RECT -98.235000  -2.300000 -98.065000  -2.130000 ;
      RECT -98.235000  -1.940000 -98.065000  -1.770000 ;
      RECT -98.235000  -1.580000 -98.065000  -1.410000 ;
      RECT -98.235000  -1.220000 -98.065000  -1.050000 ;
      RECT -98.235000  -0.860000 -98.065000  -0.690000 ;
      RECT -98.235000  -0.500000 -98.065000  -0.330000 ;
      RECT -98.235000  -0.140000 -98.065000   0.030000 ;
      RECT -98.235000   0.220000 -98.065000   0.390000 ;
      RECT -98.235000   0.580000 -98.065000   0.750000 ;
      RECT -98.235000   0.940000 -98.065000   1.110000 ;
      RECT -98.235000   1.300000 -98.065000   1.470000 ;
      RECT -98.235000   1.660000 -98.065000   1.830000 ;
      RECT -98.235000   2.020000 -98.065000   2.190000 ;
      RECT -98.235000   2.380000 -98.065000   2.550000 ;
      RECT -98.235000   2.740000 -98.065000   2.910000 ;
      RECT -98.235000   3.100000 -98.065000   3.270000 ;
      RECT -98.235000   3.460000 -98.065000   3.630000 ;
      RECT -98.235000   3.820000 -98.065000   3.990000 ;
      RECT -98.235000   4.180000 -98.065000   4.350000 ;
      RECT -98.235000   4.540000 -98.065000   4.710000 ;
      RECT -98.235000   4.900000 -98.065000   5.070000 ;
      RECT -98.235000   5.260000 -98.065000   5.430000 ;
      RECT -98.235000   5.620000 -98.065000   5.790000 ;
      RECT -98.235000   5.980000 -98.065000   6.150000 ;
      RECT -98.235000   6.340000 -98.065000   6.510000 ;
      RECT -98.235000   6.700000 -98.065000   6.870000 ;
      RECT -98.235000   7.060000 -98.065000   7.230000 ;
      RECT -98.235000   7.420000 -98.065000   7.590000 ;
      RECT -98.235000   7.780000 -98.065000   7.950000 ;
      RECT -98.235000   8.140000 -98.065000   8.310000 ;
      RECT -98.235000   8.500000 -98.065000   8.670000 ;
      RECT -98.235000   8.860000 -98.065000   9.030000 ;
      RECT -98.235000   9.220000 -98.065000   9.390000 ;
      RECT -98.235000   9.580000 -98.065000   9.750000 ;
      RECT -98.235000   9.940000 -98.065000  10.110000 ;
      RECT -98.235000  10.300000 -98.065000  10.470000 ;
      RECT -98.235000  10.660000 -98.065000  10.830000 ;
      RECT -98.235000  11.020000 -98.065000  11.190000 ;
      RECT -98.235000  11.380000 -98.065000  11.550000 ;
      RECT -98.235000  11.740000 -98.065000  11.910000 ;
      RECT -98.235000  12.100000 -98.065000  12.270000 ;
      RECT -98.235000  12.460000 -98.065000  12.630000 ;
      RECT -98.235000  12.820000 -98.065000  12.990000 ;
      RECT -98.235000  13.180000 -98.065000  13.350000 ;
      RECT -98.235000  13.540000 -98.065000  13.710000 ;
      RECT -98.235000  13.900000 -98.065000  14.070000 ;
      RECT -98.235000  14.260000 -98.065000  14.430000 ;
      RECT -98.235000  14.620000 -98.065000  14.790000 ;
      RECT -98.235000  14.980000 -98.065000  15.150000 ;
      RECT -98.235000  15.340000 -98.065000  15.510000 ;
      RECT -98.235000  15.700000 -98.065000  15.870000 ;
      RECT -98.235000  16.060000 -98.065000  16.230000 ;
      RECT -98.235000  16.420000 -98.065000  16.590000 ;
      RECT -98.235000  16.780000 -98.065000  16.950000 ;
      RECT -98.235000  17.140000 -98.065000  17.310000 ;
      RECT -98.235000  17.500000 -98.065000  17.670000 ;
      RECT -98.235000  17.860000 -98.065000  18.030000 ;
      RECT -98.235000  18.220000 -98.065000  18.390000 ;
      RECT -98.235000  18.580000 -98.065000  18.750000 ;
      RECT -98.235000  18.940000 -98.065000  19.110000 ;
      RECT -98.235000  19.300000 -98.065000  19.470000 ;
      RECT -98.235000  19.660000 -98.065000  19.830000 ;
      RECT -98.235000  20.020000 -98.065000  20.190000 ;
      RECT -98.235000  20.380000 -98.065000  20.550000 ;
      RECT -98.235000  20.740000 -98.065000  20.910000 ;
      RECT -98.235000  21.100000 -98.065000  21.270000 ;
      RECT -98.235000  21.460000 -98.065000  21.630000 ;
      RECT -98.235000  21.820000 -98.065000  21.990000 ;
      RECT -98.235000  22.180000 -98.065000  22.350000 ;
      RECT -98.235000  22.540000 -98.065000  22.710000 ;
      RECT -98.235000  22.900000 -98.065000  23.070000 ;
      RECT -98.235000  23.260000 -98.065000  23.430000 ;
      RECT -98.235000  23.620000 -98.065000  23.790000 ;
      RECT -98.235000  23.980000 -98.065000  24.150000 ;
      RECT -98.235000  24.340000 -98.065000  24.510000 ;
      RECT -98.235000  24.700000 -98.065000  24.870000 ;
      RECT -98.235000  25.060000 -98.065000  25.230000 ;
      RECT -98.235000  25.420000 -98.065000  25.590000 ;
      RECT -98.235000  25.780000 -98.065000  25.950000 ;
      RECT -98.235000  26.140000 -98.065000  26.310000 ;
      RECT -98.235000  26.500000 -98.065000  26.670000 ;
      RECT -98.235000  26.860000 -98.065000  27.030000 ;
      RECT -98.235000  27.220000 -98.065000  27.390000 ;
      RECT -98.235000  27.580000 -98.065000  27.750000 ;
      RECT -98.235000  27.940000 -98.065000  28.110000 ;
      RECT -98.235000  28.300000 -98.065000  28.470000 ;
      RECT -98.235000  28.660000 -98.065000  28.830000 ;
      RECT -98.235000  29.020000 -98.065000  29.190000 ;
      RECT -98.235000  29.380000 -98.065000  29.550000 ;
      RECT -98.235000  29.740000 -98.065000  29.910000 ;
      RECT -98.235000  30.100000 -98.065000  30.270000 ;
      RECT -98.235000  30.460000 -98.065000  30.630000 ;
      RECT -98.235000  30.820000 -98.065000  30.990000 ;
      RECT -98.235000  31.180000 -98.065000  31.350000 ;
      RECT -98.235000  31.540000 -98.065000  31.710000 ;
      RECT -98.235000  31.900000 -98.065000  32.070000 ;
      RECT -98.235000  32.260000 -98.065000  32.430000 ;
      RECT -98.235000  32.620000 -98.065000  32.790000 ;
      RECT -98.235000  32.980000 -98.065000  33.150000 ;
      RECT -98.235000  33.340000 -98.065000  33.510000 ;
      RECT -98.235000  33.700000 -98.065000  33.870000 ;
      RECT -98.235000  34.060000 -98.065000  34.230000 ;
      RECT -98.235000  34.420000 -98.065000  34.590000 ;
      RECT -98.235000  34.780000 -98.065000  34.950000 ;
      RECT -98.235000  35.140000 -98.065000  35.310000 ;
      RECT -98.235000  35.500000 -98.065000  35.670000 ;
      RECT -98.235000  35.860000 -98.065000  36.030000 ;
      RECT -98.235000  36.220000 -98.065000  36.390000 ;
      RECT -98.235000  36.580000 -98.065000  36.750000 ;
      RECT -98.235000  36.940000 -98.065000  37.110000 ;
      RECT -98.235000  37.300000 -98.065000  37.470000 ;
      RECT -98.235000  37.660000 -98.065000  37.830000 ;
      RECT -98.235000  38.020000 -98.065000  38.190000 ;
      RECT -98.235000  38.380000 -98.065000  38.550000 ;
      RECT -98.235000  38.740000 -98.065000  38.910000 ;
      RECT -98.235000  39.100000 -98.065000  39.270000 ;
      RECT -98.235000  39.460000 -98.065000  39.630000 ;
      RECT -98.235000  39.820000 -98.065000  39.990000 ;
      RECT -98.235000  40.180000 -98.065000  40.350000 ;
      RECT -98.235000  40.540000 -98.065000  40.710000 ;
      RECT -98.235000  40.900000 -98.065000  41.070000 ;
      RECT -98.235000  41.260000 -98.065000  41.430000 ;
      RECT -98.235000  41.620000 -98.065000  41.790000 ;
      RECT -98.235000  41.980000 -98.065000  42.150000 ;
      RECT -98.235000  42.340000 -98.065000  42.510000 ;
      RECT -98.235000  42.700000 -98.065000  42.870000 ;
      RECT -98.235000  43.060000 -98.065000  43.230000 ;
      RECT -98.235000  43.420000 -98.065000  43.590000 ;
      RECT -98.235000  43.780000 -98.065000  43.950000 ;
      RECT -98.235000  44.140000 -98.065000  44.310000 ;
      RECT -98.235000  44.500000 -98.065000  44.670000 ;
      RECT -98.235000  44.860000 -98.065000  45.030000 ;
      RECT -98.235000  45.220000 -98.065000  45.390000 ;
      RECT -98.235000  45.580000 -98.065000  45.750000 ;
      RECT -98.235000  45.940000 -98.065000  46.110000 ;
      RECT -98.235000  46.300000 -98.065000  46.470000 ;
      RECT -98.235000  46.660000 -98.065000  46.830000 ;
      RECT -98.235000  47.020000 -98.065000  47.190000 ;
      RECT -98.235000  47.380000 -98.065000  47.550000 ;
      RECT -98.235000  47.740000 -98.065000  47.910000 ;
      RECT -98.235000  48.100000 -98.065000  48.270000 ;
      RECT -98.235000  48.460000 -98.065000  48.630000 ;
      RECT -98.235000  48.820000 -98.065000  48.990000 ;
      RECT -98.235000  49.180000 -98.065000  49.350000 ;
      RECT -98.235000  49.540000 -98.065000  49.710000 ;
      RECT -98.235000  49.900000 -98.065000  50.070000 ;
      RECT -98.235000  50.260000 -98.065000  50.430000 ;
      RECT -98.235000  50.620000 -98.065000  50.790000 ;
      RECT -98.235000  50.980000 -98.065000  51.150000 ;
      RECT -98.235000  51.340000 -98.065000  51.510000 ;
      RECT -98.235000  51.700000 -98.065000  51.870000 ;
      RECT -98.235000  52.060000 -98.065000  52.230000 ;
      RECT -98.235000  52.420000 -98.065000  52.590000 ;
      RECT -98.235000  52.780000 -98.065000  52.950000 ;
      RECT -98.235000  53.140000 -98.065000  53.310000 ;
      RECT -98.235000  53.500000 -98.065000  53.670000 ;
      RECT -98.235000  53.860000 -98.065000  54.030000 ;
      RECT -98.235000  54.220000 -98.065000  54.390000 ;
      RECT -98.235000  54.580000 -98.065000  54.750000 ;
      RECT -98.235000  54.940000 -98.065000  55.110000 ;
      RECT -98.235000  55.300000 -98.065000  55.470000 ;
      RECT -98.235000  55.660000 -98.065000  55.830000 ;
      RECT -98.235000  56.020000 -98.065000  56.190000 ;
      RECT -98.235000  56.380000 -98.065000  56.550000 ;
      RECT -98.235000  56.740000 -98.065000  56.910000 ;
      RECT -98.235000  57.100000 -98.065000  57.270000 ;
      RECT -98.235000  57.460000 -98.065000  57.630000 ;
      RECT -98.235000  57.820000 -98.065000  57.990000 ;
      RECT -98.235000  58.180000 -98.065000  58.350000 ;
      RECT -98.235000  58.540000 -98.065000  58.710000 ;
      RECT -98.235000  58.900000 -98.065000  59.070000 ;
      RECT -98.235000  59.260000 -98.065000  59.430000 ;
      RECT -98.235000  59.620000 -98.065000  59.790000 ;
      RECT -98.235000  59.980000 -98.065000  60.150000 ;
      RECT -98.235000  60.340000 -98.065000  60.510000 ;
      RECT -98.235000  60.700000 -98.065000  60.870000 ;
      RECT -98.235000  61.060000 -98.065000  61.230000 ;
      RECT -98.235000  61.420000 -98.065000  61.590000 ;
      RECT -98.235000  61.780000 -98.065000  61.950000 ;
      RECT -98.235000  62.140000 -98.065000  62.310000 ;
      RECT -98.235000  62.500000 -98.065000  62.670000 ;
      RECT -98.235000  62.860000 -98.065000  63.030000 ;
      RECT -98.235000  63.220000 -98.065000  63.390000 ;
      RECT -98.235000  63.580000 -98.065000  63.750000 ;
      RECT -98.235000  63.940000 -98.065000  64.110000 ;
      RECT -98.235000  64.300000 -98.065000  64.470000 ;
      RECT -98.235000  64.660000 -98.065000  64.830000 ;
      RECT -98.235000  65.020000 -98.065000  65.190000 ;
      RECT -98.235000  65.380000 -98.065000  65.550000 ;
      RECT -98.235000  65.740000 -98.065000  65.910000 ;
      RECT -98.235000  66.100000 -98.065000  66.270000 ;
      RECT -98.235000  66.460000 -98.065000  66.630000 ;
      RECT -98.235000  66.820000 -98.065000  66.990000 ;
      RECT -98.235000  67.180000 -98.065000  67.350000 ;
      RECT -98.235000  67.540000 -98.065000  67.710000 ;
      RECT -98.235000  67.900000 -98.065000  68.070000 ;
      RECT -98.235000  68.260000 -98.065000  68.430000 ;
      RECT -98.235000  68.620000 -98.065000  68.790000 ;
      RECT -98.235000  68.980000 -98.065000  69.150000 ;
      RECT -98.235000  69.340000 -98.065000  69.510000 ;
      RECT -98.235000  69.700000 -98.065000  69.870000 ;
      RECT -98.235000  70.060000 -98.065000  70.230000 ;
      RECT -98.235000  70.420000 -98.065000  70.590000 ;
      RECT -98.235000  70.780000 -98.065000  70.950000 ;
      RECT -98.235000  71.140000 -98.065000  71.310000 ;
      RECT -98.235000  71.500000 -98.065000  71.670000 ;
      RECT -98.235000  71.860000 -98.065000  72.030000 ;
      RECT -98.235000  72.220000 -98.065000  72.390000 ;
      RECT -98.235000  72.580000 -98.065000  72.750000 ;
      RECT -98.235000  72.940000 -98.065000  73.110000 ;
      RECT -98.235000  73.300000 -98.065000  73.470000 ;
      RECT -98.235000  73.660000 -98.065000  73.830000 ;
      RECT -98.235000  74.020000 -98.065000  74.190000 ;
      RECT -98.235000  74.380000 -98.065000  74.550000 ;
      RECT -98.235000  74.740000 -98.065000  74.910000 ;
      RECT -98.235000  75.100000 -98.065000  75.270000 ;
      RECT -98.235000  75.460000 -98.065000  75.630000 ;
      RECT -98.235000  75.820000 -98.065000  75.990000 ;
      RECT -98.235000  76.180000 -98.065000  76.350000 ;
      RECT -98.235000  76.540000 -98.065000  76.710000 ;
      RECT -98.235000  76.900000 -98.065000  77.070000 ;
      RECT -98.235000  77.260000 -98.065000  77.430000 ;
      RECT -98.235000  77.620000 -98.065000  77.790000 ;
      RECT -98.235000  77.980000 -98.065000  78.150000 ;
      RECT -98.235000  78.340000 -98.065000  78.510000 ;
      RECT -98.235000  78.700000 -98.065000  78.870000 ;
      RECT -98.235000  79.060000 -98.065000  79.230000 ;
      RECT -98.235000  79.420000 -98.065000  79.590000 ;
      RECT -98.235000  79.780000 -98.065000  79.950000 ;
      RECT -98.235000  80.140000 -98.065000  80.310000 ;
      RECT -98.235000  80.500000 -98.065000  80.670000 ;
      RECT -98.235000  80.860000 -98.065000  81.030000 ;
      RECT -98.235000  81.220000 -98.065000  81.390000 ;
      RECT -98.235000  81.580000 -98.065000  81.750000 ;
      RECT -98.235000  81.940000 -98.065000  82.110000 ;
      RECT -98.235000  82.300000 -98.065000  82.470000 ;
      RECT -98.235000  82.660000 -98.065000  82.830000 ;
      RECT -98.235000  83.020000 -98.065000  83.190000 ;
      RECT -98.235000  83.380000 -98.065000  83.550000 ;
      RECT -98.235000  83.740000 -98.065000  83.910000 ;
      RECT -98.235000  84.100000 -98.065000  84.270000 ;
      RECT -98.235000  84.460000 -98.065000  84.630000 ;
      RECT -98.235000  84.820000 -98.065000  84.990000 ;
      RECT -98.235000  85.180000 -98.065000  85.350000 ;
      RECT -98.235000  85.540000 -98.065000  85.710000 ;
      RECT -98.235000  85.900000 -98.065000  86.070000 ;
      RECT -98.235000  86.260000 -98.065000  86.430000 ;
      RECT -98.235000  86.620000 -98.065000  86.790000 ;
      RECT -98.235000  86.980000 -98.065000  87.150000 ;
      RECT -98.235000  87.340000 -98.065000  87.510000 ;
      RECT -98.235000  87.700000 -98.065000  87.870000 ;
      RECT -98.235000  88.060000 -98.065000  88.230000 ;
      RECT -98.235000  88.420000 -98.065000  88.590000 ;
      RECT -98.235000  88.780000 -98.065000  88.950000 ;
      RECT -98.235000  89.140000 -98.065000  89.310000 ;
      RECT -98.235000  89.500000 -98.065000  89.670000 ;
      RECT -98.235000  89.860000 -98.065000  90.030000 ;
      RECT -98.235000  90.220000 -98.065000  90.390000 ;
      RECT -98.235000  90.580000 -98.065000  90.750000 ;
      RECT -98.235000  90.940000 -98.065000  91.110000 ;
      RECT -98.235000  91.300000 -98.065000  91.470000 ;
      RECT -98.235000  91.660000 -98.065000  91.830000 ;
      RECT -98.235000  92.020000 -98.065000  92.190000 ;
      RECT -98.235000  92.380000 -98.065000  92.550000 ;
      RECT -98.235000  92.740000 -98.065000  92.910000 ;
      RECT -98.235000  93.100000 -98.065000  93.270000 ;
      RECT -98.235000  93.460000 -98.065000  93.630000 ;
      RECT -98.235000  93.820000 -98.065000  93.990000 ;
      RECT -98.235000  94.180000 -98.065000  94.350000 ;
      RECT -98.235000  94.540000 -98.065000  94.710000 ;
      RECT -98.235000  94.900000 -98.065000  95.070000 ;
      RECT -98.235000  95.260000 -98.065000  95.430000 ;
      RECT -98.235000  95.620000 -98.065000  95.790000 ;
      RECT -98.235000  95.980000 -98.065000  96.150000 ;
      RECT -98.235000  96.340000 -98.065000  96.510000 ;
      RECT -98.235000  96.700000 -98.065000  96.870000 ;
      RECT -98.235000  97.060000 -98.065000  97.230000 ;
      RECT -98.235000  97.420000 -98.065000  97.590000 ;
      RECT -98.235000  97.780000 -98.065000  97.950000 ;
      RECT -98.235000  98.140000 -98.065000  98.310000 ;
      RECT -98.235000  98.500000 -98.065000  98.670000 ;
      RECT -98.235000  98.860000 -98.065000  99.030000 ;
      RECT -98.235000  99.220000 -98.065000  99.390000 ;
      RECT -98.235000  99.580000 -98.065000  99.750000 ;
      RECT -98.235000  99.940000 -98.065000 100.110000 ;
      RECT -98.235000 100.300000 -98.065000 100.470000 ;
      RECT -98.235000 100.660000 -98.065000 100.830000 ;
      RECT -98.235000 101.020000 -98.065000 101.190000 ;
      RECT -98.235000 101.380000 -98.065000 101.550000 ;
      RECT -98.235000 101.740000 -98.065000 101.910000 ;
      RECT -98.235000 102.100000 -98.065000 102.270000 ;
      RECT -98.235000 102.460000 -98.065000 102.630000 ;
      RECT -98.235000 102.820000 -98.065000 102.990000 ;
      RECT -98.235000 103.180000 -98.065000 103.350000 ;
      RECT -98.235000 103.540000 -98.065000 103.710000 ;
      RECT -98.235000 103.900000 -98.065000 104.070000 ;
      RECT -98.235000 104.260000 -98.065000 104.430000 ;
      RECT -98.235000 104.620000 -98.065000 104.790000 ;
      RECT -98.235000 104.980000 -98.065000 105.150000 ;
      RECT -98.235000 105.340000 -98.065000 105.510000 ;
      RECT -98.235000 105.700000 -98.065000 105.870000 ;
      RECT -98.235000 106.060000 -98.065000 106.230000 ;
      RECT -98.235000 106.420000 -98.065000 106.590000 ;
      RECT -98.235000 106.780000 -98.065000 106.950000 ;
      RECT -98.235000 107.140000 -98.065000 107.310000 ;
      RECT -98.235000 107.500000 -98.065000 107.670000 ;
      RECT -98.235000 107.860000 -98.065000 108.030000 ;
      RECT -98.235000 108.220000 -98.065000 108.390000 ;
      RECT -98.235000 108.580000 -98.065000 108.750000 ;
      RECT -98.235000 108.940000 -98.065000 109.110000 ;
      RECT -98.235000 109.300000 -98.065000 109.470000 ;
      RECT -98.235000 109.660000 -98.065000 109.830000 ;
      RECT -98.235000 110.020000 -98.065000 110.190000 ;
      RECT -98.235000 110.380000 -98.065000 110.550000 ;
      RECT -98.235000 110.740000 -98.065000 110.910000 ;
      RECT -98.235000 111.100000 -98.065000 111.270000 ;
      RECT -98.235000 111.460000 -98.065000 111.630000 ;
      RECT -98.235000 111.820000 -98.065000 111.990000 ;
      RECT -98.235000 112.180000 -98.065000 112.350000 ;
      RECT -98.235000 112.540000 -98.065000 112.710000 ;
      RECT -98.235000 112.900000 -98.065000 113.070000 ;
      RECT -98.235000 113.260000 -98.065000 113.430000 ;
      RECT -98.235000 113.620000 -98.065000 113.790000 ;
      RECT -98.235000 113.980000 -98.065000 114.150000 ;
      RECT -98.235000 114.340000 -98.065000 114.510000 ;
      RECT -98.235000 114.700000 -98.065000 114.870000 ;
      RECT -98.235000 115.060000 -98.065000 115.230000 ;
      RECT -98.235000 115.420000 -98.065000 115.590000 ;
      RECT -98.235000 115.780000 -98.065000 115.950000 ;
      RECT -98.235000 116.140000 -98.065000 116.310000 ;
      RECT -98.235000 116.500000 -98.065000 116.670000 ;
      RECT -98.235000 116.860000 -98.065000 117.030000 ;
      RECT -98.235000 117.220000 -98.065000 117.390000 ;
      RECT -98.235000 117.580000 -98.065000 117.750000 ;
      RECT -98.235000 117.940000 -98.065000 118.110000 ;
      RECT -98.235000 118.300000 -98.065000 118.470000 ;
      RECT -98.235000 118.660000 -98.065000 118.830000 ;
      RECT -98.235000 119.020000 -98.065000 119.190000 ;
      RECT -98.235000 119.380000 -98.065000 119.550000 ;
      RECT -98.235000 119.740000 -98.065000 119.910000 ;
      RECT -98.235000 120.100000 -98.065000 120.270000 ;
      RECT -98.235000 120.460000 -98.065000 120.630000 ;
      RECT -98.235000 120.820000 -98.065000 120.990000 ;
      RECT -98.235000 121.180000 -98.065000 121.350000 ;
      RECT -98.235000 121.540000 -98.065000 121.710000 ;
      RECT -98.235000 121.900000 -98.065000 122.070000 ;
      RECT -98.235000 122.260000 -98.065000 122.430000 ;
      RECT -98.235000 122.620000 -98.065000 122.790000 ;
      RECT -98.235000 122.980000 -98.065000 123.150000 ;
      RECT -98.235000 123.340000 -98.065000 123.510000 ;
      RECT -98.235000 123.700000 -98.065000 123.870000 ;
      RECT -98.235000 124.060000 -98.065000 124.230000 ;
      RECT -98.235000 124.420000 -98.065000 124.590000 ;
      RECT -98.235000 124.780000 -98.065000 124.950000 ;
      RECT -98.235000 125.140000 -98.065000 125.310000 ;
      RECT -98.235000 125.500000 -98.065000 125.670000 ;
      RECT -98.235000 125.860000 -98.065000 126.030000 ;
      RECT -98.235000 126.220000 -98.065000 126.390000 ;
      RECT -98.235000 126.580000 -98.065000 126.750000 ;
      RECT -98.235000 126.940000 -98.065000 127.110000 ;
      RECT -98.235000 127.300000 -98.065000 127.470000 ;
      RECT -98.235000 127.660000 -98.065000 127.830000 ;
      RECT -98.235000 128.020000 -98.065000 128.190000 ;
      RECT -98.235000 128.380000 -98.065000 128.550000 ;
      RECT -98.235000 128.740000 -98.065000 128.910000 ;
      RECT -98.235000 129.100000 -98.065000 129.270000 ;
      RECT -98.235000 129.460000 -98.065000 129.630000 ;
      RECT -98.235000 129.820000 -98.065000 129.990000 ;
      RECT -98.235000 130.180000 -98.065000 130.350000 ;
      RECT -98.235000 130.540000 -98.065000 130.710000 ;
      RECT -98.235000 130.900000 -98.065000 131.070000 ;
      RECT -98.235000 131.260000 -98.065000 131.430000 ;
      RECT -98.235000 131.620000 -98.065000 131.790000 ;
      RECT -98.235000 131.980000 -98.065000 132.150000 ;
      RECT -98.235000 132.340000 -98.065000 132.510000 ;
      RECT -98.235000 132.700000 -98.065000 132.870000 ;
      RECT -98.235000 133.060000 -98.065000 133.230000 ;
      RECT -98.235000 133.420000 -98.065000 133.590000 ;
      RECT -98.235000 133.780000 -98.065000 133.950000 ;
      RECT -98.235000 134.140000 -98.065000 134.310000 ;
      RECT -98.235000 134.500000 -98.065000 134.670000 ;
      RECT -98.235000 134.860000 -98.065000 135.030000 ;
      RECT -98.235000 135.220000 -98.065000 135.390000 ;
      RECT -98.235000 135.580000 -98.065000 135.750000 ;
      RECT -98.235000 135.940000 -98.065000 136.110000 ;
      RECT -98.235000 136.300000 -98.065000 136.470000 ;
      RECT -98.235000 136.660000 -98.065000 136.830000 ;
      RECT -98.235000 137.020000 -98.065000 137.190000 ;
      RECT -98.235000 137.380000 -98.065000 137.550000 ;
      RECT -98.235000 137.740000 -98.065000 137.910000 ;
      RECT -98.235000 138.100000 -98.065000 138.270000 ;
      RECT -98.235000 138.460000 -98.065000 138.630000 ;
      RECT -98.235000 138.820000 -98.065000 138.990000 ;
      RECT -98.235000 139.180000 -98.065000 139.350000 ;
      RECT -98.235000 139.540000 -98.065000 139.710000 ;
      RECT -98.235000 139.905000 -98.065000 140.075000 ;
      RECT -98.235000 140.270000 -98.065000 140.440000 ;
      RECT -98.235000 140.635000 -98.065000 140.805000 ;
      RECT -98.235000 141.000000 -98.065000 141.170000 ;
      RECT -98.235000 141.365000 -98.065000 141.535000 ;
      RECT -98.235000 141.730000 -98.065000 141.900000 ;
      RECT -98.235000 142.095000 -98.065000 142.265000 ;
      RECT -98.235000 142.460000 -98.065000 142.630000 ;
      RECT -98.235000 142.825000 -98.065000 142.995000 ;
      RECT -98.235000 143.190000 -98.065000 143.360000 ;
      RECT -98.235000 143.555000 -98.065000 143.725000 ;
      RECT -98.235000 143.920000 -98.065000 144.090000 ;
      RECT -98.235000 144.285000 -98.065000 144.455000 ;
      RECT -98.235000 144.650000 -98.065000 144.820000 ;
      RECT -98.235000 145.015000 -98.065000 145.185000 ;
      RECT -98.235000 145.380000 -98.065000 145.550000 ;
      RECT -98.235000 145.745000 -98.065000 145.915000 ;
      RECT -98.235000 146.110000 -98.065000 146.280000 ;
      RECT -98.235000 146.475000 -98.065000 146.645000 ;
      RECT -98.235000 146.840000 -98.065000 147.010000 ;
      RECT -98.235000 147.205000 -98.065000 147.375000 ;
      RECT -98.235000 147.570000 -98.065000 147.740000 ;
      RECT -98.235000 147.935000 -98.065000 148.105000 ;
      RECT -98.235000 148.300000 -98.065000 148.470000 ;
      RECT -98.235000 148.665000 -98.065000 148.835000 ;
      RECT -98.235000 149.030000 -98.065000 149.200000 ;
      RECT -98.235000 149.395000 -98.065000 149.565000 ;
      RECT -98.235000 149.760000 -98.065000 149.930000 ;
      RECT -98.235000 150.125000 -98.065000 150.295000 ;
      RECT -98.235000 150.490000 -98.065000 150.660000 ;
      RECT -98.235000 150.855000 -98.065000 151.025000 ;
      RECT -98.235000 151.220000 -98.065000 151.390000 ;
      RECT -98.235000 151.585000 -98.065000 151.755000 ;
      RECT -98.235000 151.950000 -98.065000 152.120000 ;
      RECT -98.235000 152.315000 -98.065000 152.485000 ;
      RECT -98.235000 152.680000 -98.065000 152.850000 ;
      RECT -98.235000 153.045000 -98.065000 153.215000 ;
      RECT -98.235000 153.410000 -98.065000 153.580000 ;
      RECT -98.235000 153.775000 -98.065000 153.945000 ;
      RECT -98.235000 154.140000 -98.065000 154.310000 ;
      RECT -98.235000 154.505000 -98.065000 154.675000 ;
      RECT -98.235000 154.870000 -98.065000 155.040000 ;
      RECT -98.235000 155.235000 -98.065000 155.405000 ;
      RECT -98.235000 155.600000 -98.065000 155.770000 ;
      RECT -98.235000 155.965000 -98.065000 156.135000 ;
      RECT -98.235000 156.330000 -98.065000 156.500000 ;
      RECT -98.150000  -8.145000 -97.980000  -7.975000 ;
      RECT -97.790000 156.415000 -97.620000 156.585000 ;
      RECT -97.785000  -8.145000 -97.615000  -7.975000 ;
      RECT -97.430000 156.415000 -97.260000 156.585000 ;
      RECT -97.420000  -8.145000 -97.250000  -7.975000 ;
      RECT -97.070000 156.415000 -96.900000 156.585000 ;
      RECT -97.055000  -8.145000 -96.885000  -7.975000 ;
      RECT -96.710000 156.415000 -96.540000 156.585000 ;
      RECT -96.690000  -8.145000 -96.520000  -7.975000 ;
      RECT -96.350000 156.415000 -96.180000 156.585000 ;
      RECT -96.325000  -8.145000 -96.155000  -7.975000 ;
      RECT -95.990000 156.415000 -95.820000 156.585000 ;
      RECT -95.960000  -8.145000 -95.790000  -7.975000 ;
      RECT -95.630000 156.415000 -95.460000 156.585000 ;
      RECT -95.595000  -8.145000 -95.425000  -7.975000 ;
      RECT -95.270000 156.415000 -95.100000 156.585000 ;
      RECT -95.230000  -8.145000 -95.060000  -7.975000 ;
      RECT -94.910000 156.415000 -94.740000 156.585000 ;
      RECT -94.865000  -8.145000 -94.695000  -7.975000 ;
      RECT -94.550000 156.415000 -94.380000 156.585000 ;
      RECT -94.500000  -8.145000 -94.330000  -7.975000 ;
      RECT -94.190000 156.415000 -94.020000 156.585000 ;
      RECT -94.135000  -8.145000 -93.965000  -7.975000 ;
      RECT -93.830000 156.415000 -93.660000 156.585000 ;
      RECT -93.770000  -8.145000 -93.600000  -7.975000 ;
      RECT -93.470000 156.415000 -93.300000 156.585000 ;
      RECT -93.405000  -8.145000 -93.235000  -7.975000 ;
      RECT -93.110000 156.415000 -92.940000 156.585000 ;
      RECT -93.040000  -8.145000 -92.870000  -7.975000 ;
      RECT -92.750000 156.415000 -92.580000 156.585000 ;
      RECT -92.675000  -8.145000 -92.505000  -7.975000 ;
      RECT -92.390000 156.415000 -92.220000 156.585000 ;
      RECT -92.310000  -8.145000 -92.140000  -7.975000 ;
      RECT -92.030000 156.415000 -91.860000 156.585000 ;
      RECT -91.945000  -8.145000 -91.775000  -7.975000 ;
      RECT -91.670000 156.415000 -91.500000 156.585000 ;
      RECT -91.580000  -8.145000 -91.410000  -7.975000 ;
      RECT -91.310000 156.415000 -91.140000 156.585000 ;
      RECT -91.215000  -8.145000 -91.045000  -7.975000 ;
      RECT -90.950000 156.415000 -90.780000 156.585000 ;
      RECT -90.850000  -8.145000 -90.680000  -7.975000 ;
      RECT -90.590000 156.415000 -90.420000 156.585000 ;
      RECT -90.485000  -8.145000 -90.315000  -7.975000 ;
      RECT -90.230000 156.415000 -90.060000 156.585000 ;
      RECT -90.120000  -8.145000 -89.950000  -7.975000 ;
      RECT -89.870000 156.415000 -89.700000 156.585000 ;
      RECT -89.755000  -8.145000 -89.585000  -7.975000 ;
      RECT -89.510000 156.415000 -89.340000 156.585000 ;
      RECT -89.390000  -8.145000 -89.220000  -7.975000 ;
      RECT -89.150000 156.415000 -88.980000 156.585000 ;
      RECT -89.025000  -8.145000 -88.855000  -7.975000 ;
      RECT -88.790000 156.415000 -88.620000 156.585000 ;
      RECT -88.660000  -8.145000 -88.490000  -7.975000 ;
      RECT -88.430000 156.415000 -88.260000 156.585000 ;
      RECT -88.295000  -8.145000 -88.125000  -7.975000 ;
      RECT -88.070000 156.415000 -87.900000 156.585000 ;
      RECT -87.930000  -8.145000 -87.760000  -7.975000 ;
      RECT -87.710000 156.415000 -87.540000 156.585000 ;
      RECT -87.565000  -8.145000 -87.395000  -7.975000 ;
      RECT -87.350000 156.415000 -87.180000 156.585000 ;
      RECT -87.200000  -8.145000 -87.030000  -7.975000 ;
      RECT -86.990000 156.415000 -86.820000 156.585000 ;
      RECT -86.835000  -8.145000 -86.665000  -7.975000 ;
      RECT -86.630000 156.415000 -86.460000 156.585000 ;
      RECT -86.470000  -8.145000 -86.300000  -7.975000 ;
      RECT -86.270000 156.415000 -86.100000 156.585000 ;
      RECT -86.105000  -8.145000 -85.935000  -7.975000 ;
      RECT -85.910000 156.415000 -85.740000 156.585000 ;
      RECT -85.740000  -8.145000 -85.570000  -7.975000 ;
      RECT -85.550000 156.415000 -85.380000 156.585000 ;
      RECT -85.375000  -8.145000 -85.205000  -7.975000 ;
      RECT -85.190000 156.415000 -85.020000 156.585000 ;
      RECT -85.010000  -8.145000 -84.840000  -7.975000 ;
      RECT -84.830000 156.415000 -84.660000 156.585000 ;
      RECT -84.645000  -8.145000 -84.475000  -7.975000 ;
      RECT -84.470000 156.415000 -84.300000 156.585000 ;
      RECT -84.280000  -8.145000 -84.110000  -7.975000 ;
      RECT -84.110000 156.415000 -83.940000 156.585000 ;
      RECT -83.915000  -8.145000 -83.745000  -7.975000 ;
      RECT -83.750000 156.415000 -83.580000 156.585000 ;
      RECT -83.550000  -8.145000 -83.380000  -7.975000 ;
      RECT -83.390000 156.415000 -83.220000 156.585000 ;
      RECT -83.185000  -8.145000 -83.015000  -7.975000 ;
      RECT -83.030000 156.415000 -82.860000 156.585000 ;
      RECT -82.820000  -8.145000 -82.650000  -7.975000 ;
      RECT -82.670000 156.415000 -82.500000 156.585000 ;
      RECT -82.455000  -8.145000 -82.285000  -7.975000 ;
      RECT -82.310000 156.415000 -82.140000 156.585000 ;
      RECT -82.090000  -8.145000 -81.920000  -7.975000 ;
      RECT -81.950000 156.415000 -81.780000 156.585000 ;
      RECT -81.725000  -8.145000 -81.555000  -7.975000 ;
      RECT -81.590000 156.415000 -81.420000 156.585000 ;
      RECT -81.360000  -8.145000 -81.190000  -7.975000 ;
      RECT -81.230000 156.415000 -81.060000 156.585000 ;
      RECT -81.000000  -8.145000 -80.830000  -7.975000 ;
      RECT -80.870000 156.415000 -80.700000 156.585000 ;
      RECT -80.640000  -8.145000 -80.470000  -7.975000 ;
      RECT -80.510000 156.415000 -80.340000 156.585000 ;
      RECT -80.280000  -8.145000 -80.110000  -7.975000 ;
      RECT -80.150000 156.415000 -79.980000 156.585000 ;
      RECT -79.920000  -8.145000 -79.750000  -7.975000 ;
      RECT -79.790000 156.415000 -79.620000 156.585000 ;
      RECT -79.560000  -8.145000 -79.390000  -7.975000 ;
      RECT -79.430000 156.415000 -79.260000 156.585000 ;
      RECT -79.200000  -8.145000 -79.030000  -7.975000 ;
      RECT -79.070000 156.415000 -78.900000 156.585000 ;
      RECT -78.840000  -8.145000 -78.670000  -7.975000 ;
      RECT -78.710000 156.415000 -78.540000 156.585000 ;
      RECT -78.480000  -8.145000 -78.310000  -7.975000 ;
      RECT -78.350000 156.415000 -78.180000 156.585000 ;
      RECT -78.120000  -8.145000 -77.950000  -7.975000 ;
      RECT -77.990000 156.415000 -77.820000 156.585000 ;
      RECT -77.760000  -8.145000 -77.590000  -7.975000 ;
      RECT -77.630000 156.415000 -77.460000 156.585000 ;
      RECT -77.400000  -8.145000 -77.230000  -7.975000 ;
      RECT -77.270000 156.415000 -77.100000 156.585000 ;
      RECT -77.040000  -8.145000 -76.870000  -7.975000 ;
      RECT -76.910000 156.415000 -76.740000 156.585000 ;
      RECT -76.680000  -8.145000 -76.510000  -7.975000 ;
      RECT -76.550000 156.415000 -76.380000 156.585000 ;
      RECT -76.320000  -8.145000 -76.150000  -7.975000 ;
      RECT -76.190000 156.415000 -76.020000 156.585000 ;
      RECT -75.960000  -8.145000 -75.790000  -7.975000 ;
      RECT -75.830000 156.415000 -75.660000 156.585000 ;
      RECT -75.600000  -8.145000 -75.430000  -7.975000 ;
      RECT -75.470000 156.415000 -75.300000 156.585000 ;
      RECT -75.240000  -8.145000 -75.070000  -7.975000 ;
      RECT -75.110000 156.415000 -74.940000 156.585000 ;
      RECT -74.880000  -8.145000 -74.710000  -7.975000 ;
      RECT -74.750000 156.415000 -74.580000 156.585000 ;
      RECT -74.520000  -8.145000 -74.350000  -7.975000 ;
      RECT -74.390000 156.415000 -74.220000 156.585000 ;
      RECT -74.160000  -8.145000 -73.990000  -7.975000 ;
      RECT -74.030000 156.415000 -73.860000 156.585000 ;
      RECT -73.800000  -8.145000 -73.630000  -7.975000 ;
      RECT -73.670000 156.415000 -73.500000 156.585000 ;
      RECT -73.440000  -8.145000 -73.270000  -7.975000 ;
      RECT -73.310000 156.415000 -73.140000 156.585000 ;
      RECT -73.080000  -8.145000 -72.910000  -7.975000 ;
      RECT -72.950000 156.415000 -72.780000 156.585000 ;
      RECT -72.720000  -8.145000 -72.550000  -7.975000 ;
      RECT -72.590000 156.415000 -72.420000 156.585000 ;
      RECT -72.360000  -8.145000 -72.190000  -7.975000 ;
      RECT -72.230000 156.415000 -72.060000 156.585000 ;
      RECT -72.000000  -8.145000 -71.830000  -7.975000 ;
      RECT -71.870000 156.415000 -71.700000 156.585000 ;
      RECT -71.640000  -8.145000 -71.470000  -7.975000 ;
      RECT -71.510000 156.415000 -71.340000 156.585000 ;
      RECT -71.280000  -8.145000 -71.110000  -7.975000 ;
      RECT -71.150000 156.415000 -70.980000 156.585000 ;
      RECT -70.920000  -8.145000 -70.750000  -7.975000 ;
      RECT -70.790000 156.415000 -70.620000 156.585000 ;
      RECT -70.560000  -8.145000 -70.390000  -7.975000 ;
      RECT -70.430000 156.415000 -70.260000 156.585000 ;
      RECT -70.200000  -8.145000 -70.030000  -7.975000 ;
      RECT -70.070000 156.415000 -69.900000 156.585000 ;
      RECT -69.840000  -8.145000 -69.670000  -7.975000 ;
      RECT -69.710000 156.415000 -69.540000 156.585000 ;
      RECT -69.480000  -8.145000 -69.310000  -7.975000 ;
      RECT -69.350000 156.415000 -69.180000 156.585000 ;
      RECT -69.120000  -8.145000 -68.950000  -7.975000 ;
      RECT -68.990000 156.415000 -68.820000 156.585000 ;
      RECT -68.760000  -8.145000 -68.590000  -7.975000 ;
      RECT -68.630000 156.415000 -68.460000 156.585000 ;
      RECT -68.400000  -8.145000 -68.230000  -7.975000 ;
      RECT -68.270000 156.415000 -68.100000 156.585000 ;
      RECT -68.040000  -8.145000 -67.870000  -7.975000 ;
      RECT -67.910000 156.415000 -67.740000 156.585000 ;
      RECT -67.680000  -8.145000 -67.510000  -7.975000 ;
      RECT -67.550000 156.415000 -67.380000 156.585000 ;
      RECT -67.320000  -8.145000 -67.150000  -7.975000 ;
      RECT -67.190000 156.415000 -67.020000 156.585000 ;
      RECT -66.960000  -8.145000 -66.790000  -7.975000 ;
      RECT -66.830000 156.415000 -66.660000 156.585000 ;
      RECT -66.600000  -8.145000 -66.430000  -7.975000 ;
      RECT -66.470000 156.415000 -66.300000 156.585000 ;
      RECT -66.240000  -8.145000 -66.070000  -7.975000 ;
      RECT -66.110000 156.415000 -65.940000 156.585000 ;
      RECT -65.880000  -8.145000 -65.710000  -7.975000 ;
      RECT -65.750000 156.415000 -65.580000 156.585000 ;
      RECT -65.520000  -8.145000 -65.350000  -7.975000 ;
      RECT -65.390000 156.415000 -65.220000 156.585000 ;
      RECT -65.160000  -8.145000 -64.990000  -7.975000 ;
      RECT -65.030000 156.415000 -64.860000 156.585000 ;
      RECT -64.800000  -8.145000 -64.630000  -7.975000 ;
      RECT -64.670000 156.415000 -64.500000 156.585000 ;
      RECT -64.440000  -8.145000 -64.270000  -7.975000 ;
      RECT -64.310000 156.415000 -64.140000 156.585000 ;
      RECT -64.080000  -8.145000 -63.910000  -7.975000 ;
      RECT -63.950000 156.415000 -63.780000 156.585000 ;
      RECT -63.720000  -8.145000 -63.550000  -7.975000 ;
      RECT -63.590000 156.415000 -63.420000 156.585000 ;
      RECT -63.360000  -8.145000 -63.190000  -7.975000 ;
      RECT -63.230000 156.415000 -63.060000 156.585000 ;
      RECT -63.000000  -8.145000 -62.830000  -7.975000 ;
      RECT -62.870000 156.415000 -62.700000 156.585000 ;
      RECT -62.640000  -8.145000 -62.470000  -7.975000 ;
      RECT -62.510000 156.415000 -62.340000 156.585000 ;
      RECT -62.280000  -8.145000 -62.110000  -7.975000 ;
      RECT -62.150000 156.415000 -61.980000 156.585000 ;
      RECT -61.920000  -8.145000 -61.750000  -7.975000 ;
      RECT -61.790000 156.415000 -61.620000 156.585000 ;
      RECT -61.560000  -8.145000 -61.390000  -7.975000 ;
      RECT -61.430000 156.415000 -61.260000 156.585000 ;
      RECT -61.200000  -8.145000 -61.030000  -7.975000 ;
      RECT -61.070000 156.415000 -60.900000 156.585000 ;
      RECT -60.840000  -8.145000 -60.670000  -7.975000 ;
      RECT -60.710000 156.415000 -60.540000 156.585000 ;
      RECT -60.480000  -8.145000 -60.310000  -7.975000 ;
      RECT -60.350000 156.415000 -60.180000 156.585000 ;
      RECT -60.120000  -8.145000 -59.950000  -7.975000 ;
      RECT -59.990000 156.415000 -59.820000 156.585000 ;
      RECT -59.760000  -8.145000 -59.590000  -7.975000 ;
      RECT -59.630000 156.415000 -59.460000 156.585000 ;
      RECT -59.400000  -8.145000 -59.230000  -7.975000 ;
      RECT -59.270000 156.415000 -59.100000 156.585000 ;
      RECT -59.040000  -8.145000 -58.870000  -7.975000 ;
      RECT -58.910000 156.415000 -58.740000 156.585000 ;
      RECT -58.680000  -8.145000 -58.510000  -7.975000 ;
      RECT -58.550000 156.415000 -58.380000 156.585000 ;
      RECT -58.320000  -8.145000 -58.150000  -7.975000 ;
      RECT -58.190000 156.415000 -58.020000 156.585000 ;
      RECT -57.960000  -8.145000 -57.790000  -7.975000 ;
      RECT -57.830000 156.415000 -57.660000 156.585000 ;
      RECT -57.600000  -8.145000 -57.430000  -7.975000 ;
      RECT -57.470000 156.415000 -57.300000 156.585000 ;
      RECT -57.240000  -8.145000 -57.070000  -7.975000 ;
      RECT -57.110000 156.415000 -56.940000 156.585000 ;
      RECT -56.880000  -8.145000 -56.710000  -7.975000 ;
      RECT -56.750000 156.415000 -56.580000 156.585000 ;
      RECT -56.520000  -8.145000 -56.350000  -7.975000 ;
      RECT -56.390000 156.415000 -56.220000 156.585000 ;
      RECT -56.160000  -8.145000 -55.990000  -7.975000 ;
      RECT -56.030000 156.415000 -55.860000 156.585000 ;
      RECT -55.800000  -8.145000 -55.630000  -7.975000 ;
      RECT -55.670000 156.415000 -55.500000 156.585000 ;
      RECT -55.440000  -8.145000 -55.270000  -7.975000 ;
      RECT -55.310000 156.415000 -55.140000 156.585000 ;
      RECT -55.080000  -8.145000 -54.910000  -7.975000 ;
      RECT -54.950000 156.415000 -54.780000 156.585000 ;
      RECT -54.720000  -8.145000 -54.550000  -7.975000 ;
      RECT -54.590000 156.415000 -54.420000 156.585000 ;
      RECT -54.360000  -8.145000 -54.190000  -7.975000 ;
      RECT -54.230000 156.415000 -54.060000 156.585000 ;
      RECT -54.000000  -8.145000 -53.830000  -7.975000 ;
      RECT -53.870000 156.415000 -53.700000 156.585000 ;
      RECT -53.640000  -8.145000 -53.470000  -7.975000 ;
      RECT -53.510000 156.415000 -53.340000 156.585000 ;
      RECT -53.280000  -8.145000 -53.110000  -7.975000 ;
      RECT -53.150000 156.415000 -52.980000 156.585000 ;
      RECT -52.920000  -8.145000 -52.750000  -7.975000 ;
      RECT -52.790000 156.415000 -52.620000 156.585000 ;
      RECT -52.560000  -8.145000 -52.390000  -7.975000 ;
      RECT -52.430000 156.415000 -52.260000 156.585000 ;
      RECT -52.200000  -8.145000 -52.030000  -7.975000 ;
      RECT -52.070000 156.415000 -51.900000 156.585000 ;
      RECT -51.840000  -8.145000 -51.670000  -7.975000 ;
      RECT -51.710000 156.415000 -51.540000 156.585000 ;
      RECT -51.480000  -8.145000 -51.310000  -7.975000 ;
      RECT -51.350000 156.415000 -51.180000 156.585000 ;
      RECT -51.120000  -8.145000 -50.950000  -7.975000 ;
      RECT -50.990000 156.415000 -50.820000 156.585000 ;
      RECT -50.760000  -8.145000 -50.590000  -7.975000 ;
      RECT -50.630000 156.415000 -50.460000 156.585000 ;
      RECT -50.400000  -8.145000 -50.230000  -7.975000 ;
      RECT -50.270000 156.415000 -50.100000 156.585000 ;
      RECT -50.040000  -8.145000 -49.870000  -7.975000 ;
      RECT -49.910000 156.415000 -49.740000 156.585000 ;
      RECT -49.680000  -8.145000 -49.510000  -7.975000 ;
      RECT -49.550000 156.415000 -49.380000 156.585000 ;
      RECT -49.320000  -8.145000 -49.150000  -7.975000 ;
      RECT -49.190000 156.415000 -49.020000 156.585000 ;
      RECT -48.960000  -8.145000 -48.790000  -7.975000 ;
      RECT -48.830000 156.415000 -48.660000 156.585000 ;
      RECT -48.600000  -8.145000 -48.430000  -7.975000 ;
      RECT -48.470000 156.415000 -48.300000 156.585000 ;
      RECT -48.240000  -8.145000 -48.070000  -7.975000 ;
      RECT -48.110000 156.415000 -47.940000 156.585000 ;
      RECT -47.880000  -8.145000 -47.710000  -7.975000 ;
      RECT -47.750000 156.415000 -47.580000 156.585000 ;
      RECT -47.520000  -8.145000 -47.350000  -7.975000 ;
      RECT -47.390000 156.415000 -47.220000 156.585000 ;
      RECT -47.160000  -8.145000 -46.990000  -7.975000 ;
      RECT -47.030000 156.415000 -46.860000 156.585000 ;
      RECT -46.800000  -8.145000 -46.630000  -7.975000 ;
      RECT -46.670000 156.415000 -46.500000 156.585000 ;
      RECT -46.440000  -8.145000 -46.270000  -7.975000 ;
      RECT -46.310000 156.415000 -46.140000 156.585000 ;
      RECT -46.080000  -8.145000 -45.910000  -7.975000 ;
      RECT -45.950000 156.415000 -45.780000 156.585000 ;
      RECT -45.720000  -8.145000 -45.550000  -7.975000 ;
      RECT -45.590000 156.415000 -45.420000 156.585000 ;
      RECT -45.360000  -8.145000 -45.190000  -7.975000 ;
      RECT -45.230000 156.415000 -45.060000 156.585000 ;
      RECT -45.000000  -8.145000 -44.830000  -7.975000 ;
      RECT -44.870000 156.415000 -44.700000 156.585000 ;
      RECT -44.640000  -8.145000 -44.470000  -7.975000 ;
      RECT -44.510000 156.415000 -44.340000 156.585000 ;
      RECT -44.280000  -8.145000 -44.110000  -7.975000 ;
      RECT -44.150000 156.415000 -43.980000 156.585000 ;
      RECT -43.920000  -8.145000 -43.750000  -7.975000 ;
      RECT -43.790000 156.415000 -43.620000 156.585000 ;
      RECT -43.560000  -8.145000 -43.390000  -7.975000 ;
      RECT -43.430000 156.415000 -43.260000 156.585000 ;
      RECT -43.200000  -8.145000 -43.030000  -7.975000 ;
      RECT -43.070000 156.415000 -42.900000 156.585000 ;
      RECT -42.840000  -8.145000 -42.670000  -7.975000 ;
      RECT -42.710000 156.415000 -42.540000 156.585000 ;
      RECT -42.480000  -8.145000 -42.310000  -7.975000 ;
      RECT -42.350000 156.415000 -42.180000 156.585000 ;
      RECT -42.120000  -8.145000 -41.950000  -7.975000 ;
      RECT -41.990000 156.415000 -41.820000 156.585000 ;
      RECT -41.760000  -8.145000 -41.590000  -7.975000 ;
      RECT -41.630000 156.415000 -41.460000 156.585000 ;
      RECT -41.400000  -8.145000 -41.230000  -7.975000 ;
      RECT -41.270000 156.415000 -41.100000 156.585000 ;
      RECT -41.040000  -8.145000 -40.870000  -7.975000 ;
      RECT -40.910000 156.415000 -40.740000 156.585000 ;
      RECT -40.680000  -8.145000 -40.510000  -7.975000 ;
      RECT -40.550000 156.415000 -40.380000 156.585000 ;
      RECT -40.320000  -8.145000 -40.150000  -7.975000 ;
      RECT -40.190000 156.415000 -40.020000 156.585000 ;
      RECT -39.960000  -8.145000 -39.790000  -7.975000 ;
      RECT -39.830000 156.415000 -39.660000 156.585000 ;
      RECT -39.600000  -8.145000 -39.430000  -7.975000 ;
      RECT -39.470000 156.415000 -39.300000 156.585000 ;
      RECT -39.240000  -8.145000 -39.070000  -7.975000 ;
      RECT -39.110000 156.415000 -38.940000 156.585000 ;
      RECT -38.880000  -8.145000 -38.710000  -7.975000 ;
      RECT -38.750000 156.415000 -38.580000 156.585000 ;
      RECT -38.520000  -8.145000 -38.350000  -7.975000 ;
      RECT -38.390000 156.415000 -38.220000 156.585000 ;
      RECT -38.160000  -8.145000 -37.990000  -7.975000 ;
      RECT -38.030000 156.415000 -37.860000 156.585000 ;
      RECT -37.800000  -8.145000 -37.630000  -7.975000 ;
      RECT -37.670000 156.415000 -37.500000 156.585000 ;
      RECT -37.440000  -8.145000 -37.270000  -7.975000 ;
      RECT -37.310000 156.415000 -37.140000 156.585000 ;
      RECT -37.080000  -8.145000 -36.910000  -7.975000 ;
      RECT -36.950000 156.415000 -36.780000 156.585000 ;
      RECT -36.720000  -8.145000 -36.550000  -7.975000 ;
      RECT -36.590000 156.415000 -36.420000 156.585000 ;
      RECT -36.360000  -8.145000 -36.190000  -7.975000 ;
      RECT -36.230000 156.415000 -36.060000 156.585000 ;
      RECT -36.000000  -8.145000 -35.830000  -7.975000 ;
      RECT -35.870000 156.415000 -35.700000 156.585000 ;
      RECT -35.640000  -8.145000 -35.470000  -7.975000 ;
      RECT -35.510000 156.415000 -35.340000 156.585000 ;
      RECT -35.280000  -8.145000 -35.110000  -7.975000 ;
      RECT -35.150000 156.415000 -34.980000 156.585000 ;
      RECT -34.920000  -8.145000 -34.750000  -7.975000 ;
      RECT -34.790000 156.415000 -34.620000 156.585000 ;
      RECT -34.560000  -8.145000 -34.390000  -7.975000 ;
      RECT -34.430000 156.415000 -34.260000 156.585000 ;
      RECT -34.200000  -8.145000 -34.030000  -7.975000 ;
      RECT -34.070000 156.415000 -33.900000 156.585000 ;
      RECT -33.840000  -8.145000 -33.670000  -7.975000 ;
      RECT -33.710000 156.415000 -33.540000 156.585000 ;
      RECT -33.480000  -8.145000 -33.310000  -7.975000 ;
      RECT -33.350000 156.415000 -33.180000 156.585000 ;
      RECT -33.120000  -8.145000 -32.950000  -7.975000 ;
      RECT -32.990000 156.415000 -32.820000 156.585000 ;
      RECT -32.760000  -8.145000 -32.590000  -7.975000 ;
      RECT -32.630000 156.415000 -32.460000 156.585000 ;
      RECT -32.400000  -8.145000 -32.230000  -7.975000 ;
      RECT -32.270000 156.415000 -32.100000 156.585000 ;
      RECT -32.040000  -8.145000 -31.870000  -7.975000 ;
      RECT -31.910000 156.415000 -31.740000 156.585000 ;
      RECT -31.680000  -8.145000 -31.510000  -7.975000 ;
      RECT -31.550000 156.415000 -31.380000 156.585000 ;
      RECT -31.320000  -8.145000 -31.150000  -7.975000 ;
      RECT -31.190000 156.415000 -31.020000 156.585000 ;
      RECT -30.960000  -8.145000 -30.790000  -7.975000 ;
      RECT -30.830000 156.415000 -30.660000 156.585000 ;
      RECT -30.600000  -8.145000 -30.430000  -7.975000 ;
      RECT -30.470000 156.415000 -30.300000 156.585000 ;
      RECT -30.240000  -8.145000 -30.070000  -7.975000 ;
      RECT -30.110000 156.415000 -29.940000 156.585000 ;
      RECT -29.880000  -8.145000 -29.710000  -7.975000 ;
      RECT -29.750000 156.415000 -29.580000 156.585000 ;
      RECT -29.520000  -8.145000 -29.350000  -7.975000 ;
      RECT -29.390000 156.415000 -29.220000 156.585000 ;
      RECT -29.160000  -8.145000 -28.990000  -7.975000 ;
      RECT -29.030000 156.415000 -28.860000 156.585000 ;
      RECT -28.800000  -8.145000 -28.630000  -7.975000 ;
      RECT -28.670000 156.415000 -28.500000 156.585000 ;
      RECT -28.440000  -8.145000 -28.270000  -7.975000 ;
      RECT -28.310000 156.415000 -28.140000 156.585000 ;
      RECT -28.080000  -8.145000 -27.910000  -7.975000 ;
      RECT -27.950000 156.415000 -27.780000 156.585000 ;
      RECT -27.720000  -8.145000 -27.550000  -7.975000 ;
      RECT -27.590000 156.415000 -27.420000 156.585000 ;
      RECT -27.360000  -8.145000 -27.190000  -7.975000 ;
      RECT -27.230000 156.415000 -27.060000 156.585000 ;
      RECT -27.000000  -8.145000 -26.830000  -7.975000 ;
      RECT -26.870000 156.415000 -26.700000 156.585000 ;
      RECT -26.640000  -8.145000 -26.470000  -7.975000 ;
      RECT -26.510000 156.415000 -26.340000 156.585000 ;
      RECT -26.280000  -8.145000 -26.110000  -7.975000 ;
      RECT -26.150000 156.415000 -25.980000 156.585000 ;
      RECT -25.920000  -8.145000 -25.750000  -7.975000 ;
      RECT -25.790000 156.415000 -25.620000 156.585000 ;
      RECT -25.560000  -8.145000 -25.390000  -7.975000 ;
      RECT -25.430000 156.415000 -25.260000 156.585000 ;
      RECT -25.200000  -8.145000 -25.030000  -7.975000 ;
      RECT -25.070000 156.415000 -24.900000 156.585000 ;
      RECT -24.840000  -8.145000 -24.670000  -7.975000 ;
      RECT -24.710000 156.415000 -24.540000 156.585000 ;
      RECT -24.480000  -8.145000 -24.310000  -7.975000 ;
      RECT -24.350000 156.415000 -24.180000 156.585000 ;
      RECT -24.120000  -8.145000 -23.950000  -7.975000 ;
      RECT -23.990000 156.415000 -23.820000 156.585000 ;
      RECT -23.760000  -8.145000 -23.590000  -7.975000 ;
      RECT -23.630000 156.415000 -23.460000 156.585000 ;
      RECT -23.400000  -8.145000 -23.230000  -7.975000 ;
      RECT -23.270000 156.415000 -23.100000 156.585000 ;
      RECT -23.040000  -8.145000 -22.870000  -7.975000 ;
      RECT -22.910000 156.415000 -22.740000 156.585000 ;
      RECT -22.680000  -8.145000 -22.510000  -7.975000 ;
      RECT -22.550000 156.415000 -22.380000 156.585000 ;
      RECT -22.320000  -8.145000 -22.150000  -7.975000 ;
      RECT -22.190000 156.415000 -22.020000 156.585000 ;
      RECT -21.960000  -8.145000 -21.790000  -7.975000 ;
      RECT -21.830000 156.415000 -21.660000 156.585000 ;
      RECT -21.600000  -8.145000 -21.430000  -7.975000 ;
      RECT -21.470000 156.415000 -21.300000 156.585000 ;
      RECT -21.240000  -8.145000 -21.070000  -7.975000 ;
      RECT -21.110000 156.415000 -20.940000 156.585000 ;
      RECT -20.880000  -8.145000 -20.710000  -7.975000 ;
      RECT -20.750000 156.415000 -20.580000 156.585000 ;
      RECT -20.520000  -8.145000 -20.350000  -7.975000 ;
      RECT -20.390000 156.415000 -20.220000 156.585000 ;
      RECT -20.160000  -8.145000 -19.990000  -7.975000 ;
      RECT -20.030000 156.415000 -19.860000 156.585000 ;
      RECT -19.800000  -8.145000 -19.630000  -7.975000 ;
      RECT -19.670000 156.415000 -19.500000 156.585000 ;
      RECT -19.440000  -8.145000 -19.270000  -7.975000 ;
      RECT -19.310000 156.415000 -19.140000 156.585000 ;
      RECT -19.080000  -8.145000 -18.910000  -7.975000 ;
      RECT -18.950000 156.415000 -18.780000 156.585000 ;
      RECT -18.720000  -8.145000 -18.550000  -7.975000 ;
      RECT -18.590000 156.415000 -18.420000 156.585000 ;
      RECT -18.360000  -8.145000 -18.190000  -7.975000 ;
      RECT -18.230000 156.415000 -18.060000 156.585000 ;
      RECT -18.000000  -8.145000 -17.830000  -7.975000 ;
      RECT -17.870000 156.415000 -17.700000 156.585000 ;
      RECT -17.640000  -8.145000 -17.470000  -7.975000 ;
      RECT -17.510000 156.415000 -17.340000 156.585000 ;
      RECT -17.280000  -8.145000 -17.110000  -7.975000 ;
      RECT -17.150000 156.415000 -16.980000 156.585000 ;
      RECT -16.920000  -8.145000 -16.750000  -7.975000 ;
      RECT -16.790000 156.415000 -16.620000 156.585000 ;
      RECT -16.560000  -8.145000 -16.390000  -7.975000 ;
      RECT -16.430000 156.415000 -16.260000 156.585000 ;
      RECT -16.200000  -8.145000 -16.030000  -7.975000 ;
      RECT -16.070000 156.415000 -15.900000 156.585000 ;
      RECT -15.840000  -8.145000 -15.670000  -7.975000 ;
      RECT -15.710000 156.415000 -15.540000 156.585000 ;
      RECT -15.480000  -8.145000 -15.310000  -7.975000 ;
      RECT -15.350000 156.415000 -15.180000 156.585000 ;
      RECT -15.120000  -8.145000 -14.950000  -7.975000 ;
      RECT -14.990000 156.415000 -14.820000 156.585000 ;
      RECT -14.760000  -8.145000 -14.590000  -7.975000 ;
      RECT -14.630000 156.415000 -14.460000 156.585000 ;
      RECT -14.400000  -8.145000 -14.230000  -7.975000 ;
      RECT -14.270000 156.415000 -14.100000 156.585000 ;
      RECT -14.040000  -8.145000 -13.870000  -7.975000 ;
      RECT -13.910000 156.415000 -13.740000 156.585000 ;
      RECT -13.680000  -8.145000 -13.510000  -7.975000 ;
      RECT -13.550000 156.415000 -13.380000 156.585000 ;
      RECT -13.320000  -8.145000 -13.150000  -7.975000 ;
      RECT -13.190000 156.415000 -13.020000 156.585000 ;
      RECT -12.960000  -8.145000 -12.790000  -7.975000 ;
      RECT -12.830000 156.415000 -12.660000 156.585000 ;
      RECT -12.600000  -8.145000 -12.430000  -7.975000 ;
      RECT -12.470000 156.415000 -12.300000 156.585000 ;
      RECT -12.240000  -8.145000 -12.070000  -7.975000 ;
      RECT -12.110000 156.415000 -11.940000 156.585000 ;
      RECT -11.880000  -8.145000 -11.710000  -7.975000 ;
      RECT -11.750000 156.415000 -11.580000 156.585000 ;
      RECT -11.520000  -8.145000 -11.350000  -7.975000 ;
      RECT -11.390000 156.415000 -11.220000 156.585000 ;
      RECT -11.160000  -8.145000 -10.990000  -7.975000 ;
      RECT -11.030000 156.415000 -10.860000 156.585000 ;
      RECT -10.800000  -8.145000 -10.630000  -7.975000 ;
      RECT -10.670000 156.415000 -10.500000 156.585000 ;
      RECT -10.440000  -8.145000 -10.270000  -7.975000 ;
      RECT -10.310000 156.415000 -10.140000 156.585000 ;
      RECT -10.080000  -8.145000  -9.910000  -7.975000 ;
      RECT  -9.950000 156.415000  -9.780000 156.585000 ;
      RECT  -9.720000  -8.145000  -9.550000  -7.975000 ;
      RECT  -9.590000 156.415000  -9.420000 156.585000 ;
      RECT  -9.360000  -8.145000  -9.190000  -7.975000 ;
      RECT  -9.230000 156.415000  -9.060000 156.585000 ;
      RECT  -9.000000  -8.145000  -8.830000  -7.975000 ;
      RECT  -8.870000 156.415000  -8.700000 156.585000 ;
      RECT  -8.640000  -8.145000  -8.470000  -7.975000 ;
      RECT  -8.510000 156.415000  -8.340000 156.585000 ;
      RECT  -8.280000  -8.145000  -8.110000  -7.975000 ;
      RECT  -8.150000 156.415000  -7.980000 156.585000 ;
      RECT  -7.920000  -8.145000  -7.750000  -7.975000 ;
      RECT  -7.790000 156.415000  -7.620000 156.585000 ;
      RECT  -7.560000  -8.145000  -7.390000  -7.975000 ;
      RECT  -7.430000 156.415000  -7.260000 156.585000 ;
      RECT  -7.200000  -8.145000  -7.030000  -7.975000 ;
      RECT  -7.070000 156.415000  -6.900000 156.585000 ;
      RECT  -6.840000  -8.145000  -6.670000  -7.975000 ;
      RECT  -6.710000 156.415000  -6.540000 156.585000 ;
      RECT  -6.480000  -8.145000  -6.310000  -7.975000 ;
      RECT  -6.350000 156.415000  -6.180000 156.585000 ;
      RECT  -6.120000  -8.145000  -5.950000  -7.975000 ;
      RECT  -5.990000 156.415000  -5.820000 156.585000 ;
      RECT  -5.760000  -8.145000  -5.590000  -7.975000 ;
      RECT  -5.630000 156.415000  -5.460000 156.585000 ;
      RECT  -5.400000  -8.145000  -5.230000  -7.975000 ;
      RECT  -5.270000 156.415000  -5.100000 156.585000 ;
      RECT  -5.040000  -8.145000  -4.870000  -7.975000 ;
      RECT  -4.910000 156.415000  -4.740000 156.585000 ;
      RECT  -4.680000  -8.145000  -4.510000  -7.975000 ;
      RECT  -4.550000 156.415000  -4.380000 156.585000 ;
      RECT  -4.320000  -8.145000  -4.150000  -7.975000 ;
      RECT  -4.190000 156.415000  -4.020000 156.585000 ;
      RECT  -3.960000  -8.145000  -3.790000  -7.975000 ;
      RECT  -3.830000 156.415000  -3.660000 156.585000 ;
      RECT  -3.600000  -8.145000  -3.430000  -7.975000 ;
      RECT  -3.470000 156.415000  -3.300000 156.585000 ;
      RECT  -3.240000  -8.145000  -3.070000  -7.975000 ;
      RECT  -3.110000 156.415000  -2.940000 156.585000 ;
      RECT  -2.880000  -8.145000  -2.710000  -7.975000 ;
      RECT  -2.750000 156.415000  -2.580000 156.585000 ;
      RECT  -2.520000  -8.145000  -2.350000  -7.975000 ;
      RECT  -2.390000 156.415000  -2.220000 156.585000 ;
      RECT  -2.245000  -6.385000  -2.075000  -6.215000 ;
      RECT  -2.245000  -5.165000  -2.075000  -4.995000 ;
      RECT  -2.245000  -3.945000  -2.075000  -3.775000 ;
      RECT  -2.245000  -2.725000  -2.075000  -2.555000 ;
      RECT  -2.245000  -1.505000  -2.075000  -1.335000 ;
      RECT  -2.245000  -0.285000  -2.075000  -0.115000 ;
      RECT  -2.245000   0.935000  -2.075000   1.105000 ;
      RECT  -2.245000   2.155000  -2.075000   2.325000 ;
      RECT  -2.245000   3.375000  -2.075000   3.545000 ;
      RECT  -2.245000   4.595000  -2.075000   4.765000 ;
      RECT  -2.245000   5.815000  -2.075000   5.985000 ;
      RECT  -2.245000   7.035000  -2.075000   7.205000 ;
      RECT  -2.245000   8.255000  -2.075000   8.425000 ;
      RECT  -2.245000   9.475000  -2.075000   9.645000 ;
      RECT  -2.245000  10.695000  -2.075000  10.865000 ;
      RECT  -2.245000  11.915000  -2.075000  12.085000 ;
      RECT  -2.245000  13.135000  -2.075000  13.305000 ;
      RECT  -2.245000  14.355000  -2.075000  14.525000 ;
      RECT  -2.245000  15.575000  -2.075000  15.745000 ;
      RECT  -2.245000  16.795000  -2.075000  16.965000 ;
      RECT  -2.245000  18.015000  -2.075000  18.185000 ;
      RECT  -2.245000  19.235000  -2.075000  19.405000 ;
      RECT  -2.245000  20.455000  -2.075000  20.625000 ;
      RECT  -2.245000  21.675000  -2.075000  21.845000 ;
      RECT  -2.245000  22.895000  -2.075000  23.065000 ;
      RECT  -2.245000  24.115000  -2.075000  24.285000 ;
      RECT  -2.245000  25.335000  -2.075000  25.505000 ;
      RECT  -2.245000  26.555000  -2.075000  26.725000 ;
      RECT  -2.245000  27.775000  -2.075000  27.945000 ;
      RECT  -2.245000  28.995000  -2.075000  29.165000 ;
      RECT  -2.245000  30.215000  -2.075000  30.385000 ;
      RECT  -2.245000  31.435000  -2.075000  31.605000 ;
      RECT  -2.245000  32.655000  -2.075000  32.825000 ;
      RECT  -2.245000  33.875000  -2.075000  34.045000 ;
      RECT  -2.245000  35.095000  -2.075000  35.265000 ;
      RECT  -2.245000  36.315000  -2.075000  36.485000 ;
      RECT  -2.245000  37.535000  -2.075000  37.705000 ;
      RECT  -2.245000  38.755000  -2.075000  38.925000 ;
      RECT  -2.245000  39.975000  -2.075000  40.145000 ;
      RECT  -2.245000  41.195000  -2.075000  41.365000 ;
      RECT  -2.245000  42.415000  -2.075000  42.585000 ;
      RECT  -2.245000  43.635000  -2.075000  43.805000 ;
      RECT  -2.245000  44.855000  -2.075000  45.025000 ;
      RECT  -2.245000  46.075000  -2.075000  46.245000 ;
      RECT  -2.245000  47.295000  -2.075000  47.465000 ;
      RECT  -2.245000  48.515000  -2.075000  48.685000 ;
      RECT  -2.245000  49.735000  -2.075000  49.905000 ;
      RECT  -2.245000  50.955000  -2.075000  51.125000 ;
      RECT  -2.245000  52.175000  -2.075000  52.345000 ;
      RECT  -2.245000  53.395000  -2.075000  53.565000 ;
      RECT  -2.245000  54.615000  -2.075000  54.785000 ;
      RECT  -2.245000  55.835000  -2.075000  56.005000 ;
      RECT  -2.245000  57.055000  -2.075000  57.225000 ;
      RECT  -2.245000  58.275000  -2.075000  58.445000 ;
      RECT  -2.245000  59.495000  -2.075000  59.665000 ;
      RECT  -2.245000  60.715000  -2.075000  60.885000 ;
      RECT  -2.245000  61.935000  -2.075000  62.105000 ;
      RECT  -2.245000  63.155000  -2.075000  63.325000 ;
      RECT  -2.245000  64.375000  -2.075000  64.545000 ;
      RECT  -2.245000  65.595000  -2.075000  65.765000 ;
      RECT  -2.245000  66.815000  -2.075000  66.985000 ;
      RECT  -2.245000  68.035000  -2.075000  68.205000 ;
      RECT  -2.245000  69.255000  -2.075000  69.425000 ;
      RECT  -2.245000  70.475000  -2.075000  70.645000 ;
      RECT  -2.245000  71.695000  -2.075000  71.865000 ;
      RECT  -2.245000  72.915000  -2.075000  73.085000 ;
      RECT  -2.245000  74.135000  -2.075000  74.305000 ;
      RECT  -2.245000  75.355000  -2.075000  75.525000 ;
      RECT  -2.245000  76.575000  -2.075000  76.745000 ;
      RECT  -2.245000  77.795000  -2.075000  77.965000 ;
      RECT  -2.245000  79.015000  -2.075000  79.185000 ;
      RECT  -2.245000  80.235000  -2.075000  80.405000 ;
      RECT  -2.245000  81.455000  -2.075000  81.625000 ;
      RECT  -2.245000  82.675000  -2.075000  82.845000 ;
      RECT  -2.245000  83.895000  -2.075000  84.065000 ;
      RECT  -2.245000  85.115000  -2.075000  85.285000 ;
      RECT  -2.245000  86.335000  -2.075000  86.505000 ;
      RECT  -2.245000  87.555000  -2.075000  87.725000 ;
      RECT  -2.245000  88.775000  -2.075000  88.945000 ;
      RECT  -2.245000  89.995000  -2.075000  90.165000 ;
      RECT  -2.245000  91.215000  -2.075000  91.385000 ;
      RECT  -2.245000  92.435000  -2.075000  92.605000 ;
      RECT  -2.245000  93.655000  -2.075000  93.825000 ;
      RECT  -2.245000  94.875000  -2.075000  95.045000 ;
      RECT  -2.245000  96.095000  -2.075000  96.265000 ;
      RECT  -2.245000  97.315000  -2.075000  97.485000 ;
      RECT  -2.245000  98.535000  -2.075000  98.705000 ;
      RECT  -2.245000  99.755000  -2.075000  99.925000 ;
      RECT  -2.245000 100.975000  -2.075000 101.145000 ;
      RECT  -2.245000 102.195000  -2.075000 102.365000 ;
      RECT  -2.245000 103.415000  -2.075000 103.585000 ;
      RECT  -2.245000 104.635000  -2.075000 104.805000 ;
      RECT  -2.245000 105.855000  -2.075000 106.025000 ;
      RECT  -2.245000 107.075000  -2.075000 107.245000 ;
      RECT  -2.245000 108.295000  -2.075000 108.465000 ;
      RECT  -2.245000 109.515000  -2.075000 109.685000 ;
      RECT  -2.245000 110.735000  -2.075000 110.905000 ;
      RECT  -2.245000 111.955000  -2.075000 112.125000 ;
      RECT  -2.245000 113.175000  -2.075000 113.345000 ;
      RECT  -2.245000 114.395000  -2.075000 114.565000 ;
      RECT  -2.245000 115.615000  -2.075000 115.785000 ;
      RECT  -2.245000 116.835000  -2.075000 117.005000 ;
      RECT  -2.245000 118.055000  -2.075000 118.225000 ;
      RECT  -2.245000 119.275000  -2.075000 119.445000 ;
      RECT  -2.245000 120.495000  -2.075000 120.665000 ;
      RECT  -2.245000 121.715000  -2.075000 121.885000 ;
      RECT  -2.245000 122.935000  -2.075000 123.105000 ;
      RECT  -2.245000 124.155000  -2.075000 124.325000 ;
      RECT  -2.245000 125.375000  -2.075000 125.545000 ;
      RECT  -2.245000 126.595000  -2.075000 126.765000 ;
      RECT  -2.245000 127.815000  -2.075000 127.985000 ;
      RECT  -2.245000 129.035000  -2.075000 129.205000 ;
      RECT  -2.245000 130.255000  -2.075000 130.425000 ;
      RECT  -2.245000 131.475000  -2.075000 131.645000 ;
      RECT  -2.245000 132.695000  -2.075000 132.865000 ;
      RECT  -2.245000 133.915000  -2.075000 134.085000 ;
      RECT  -2.245000 135.135000  -2.075000 135.305000 ;
      RECT  -2.245000 136.355000  -2.075000 136.525000 ;
      RECT  -2.245000 137.575000  -2.075000 137.745000 ;
      RECT  -2.245000 138.795000  -2.075000 138.965000 ;
      RECT  -2.245000 140.015000  -2.075000 140.185000 ;
      RECT  -2.245000 141.235000  -2.075000 141.405000 ;
      RECT  -2.245000 142.455000  -2.075000 142.625000 ;
      RECT  -2.245000 143.675000  -2.075000 143.845000 ;
      RECT  -2.245000 144.895000  -2.075000 145.065000 ;
      RECT  -2.245000 146.115000  -2.075000 146.285000 ;
      RECT  -2.245000 147.335000  -2.075000 147.505000 ;
      RECT  -2.245000 148.555000  -2.075000 148.725000 ;
      RECT  -2.245000 149.775000  -2.075000 149.945000 ;
      RECT  -2.245000 150.995000  -2.075000 151.165000 ;
      RECT  -2.245000 152.215000  -2.075000 152.385000 ;
      RECT  -2.245000 153.435000  -2.075000 153.605000 ;
      RECT  -2.245000 154.655000  -2.075000 154.825000 ;
      RECT  -2.160000  -8.145000  -1.990000  -7.975000 ;
      RECT  -2.030000 156.415000  -1.860000 156.585000 ;
      RECT  -1.800000  -8.145000  -1.630000  -7.975000 ;
      RECT  -1.765000  -6.385000  -1.595000  -6.215000 ;
      RECT  -1.765000  -5.165000  -1.595000  -4.995000 ;
      RECT  -1.765000  -3.945000  -1.595000  -3.775000 ;
      RECT  -1.765000  -2.725000  -1.595000  -2.555000 ;
      RECT  -1.765000  -1.505000  -1.595000  -1.335000 ;
      RECT  -1.765000  -0.285000  -1.595000  -0.115000 ;
      RECT  -1.765000   0.935000  -1.595000   1.105000 ;
      RECT  -1.765000   2.155000  -1.595000   2.325000 ;
      RECT  -1.765000   3.375000  -1.595000   3.545000 ;
      RECT  -1.765000   4.595000  -1.595000   4.765000 ;
      RECT  -1.765000   5.815000  -1.595000   5.985000 ;
      RECT  -1.765000   7.035000  -1.595000   7.205000 ;
      RECT  -1.765000   8.255000  -1.595000   8.425000 ;
      RECT  -1.765000   9.475000  -1.595000   9.645000 ;
      RECT  -1.765000  10.695000  -1.595000  10.865000 ;
      RECT  -1.765000  11.915000  -1.595000  12.085000 ;
      RECT  -1.765000  13.135000  -1.595000  13.305000 ;
      RECT  -1.765000  14.355000  -1.595000  14.525000 ;
      RECT  -1.765000  15.575000  -1.595000  15.745000 ;
      RECT  -1.765000  16.795000  -1.595000  16.965000 ;
      RECT  -1.765000  18.015000  -1.595000  18.185000 ;
      RECT  -1.765000  19.235000  -1.595000  19.405000 ;
      RECT  -1.765000  20.455000  -1.595000  20.625000 ;
      RECT  -1.765000  21.675000  -1.595000  21.845000 ;
      RECT  -1.765000  22.895000  -1.595000  23.065000 ;
      RECT  -1.765000  24.115000  -1.595000  24.285000 ;
      RECT  -1.765000  25.335000  -1.595000  25.505000 ;
      RECT  -1.765000  26.555000  -1.595000  26.725000 ;
      RECT  -1.765000  27.775000  -1.595000  27.945000 ;
      RECT  -1.765000  28.995000  -1.595000  29.165000 ;
      RECT  -1.765000  30.215000  -1.595000  30.385000 ;
      RECT  -1.765000  31.435000  -1.595000  31.605000 ;
      RECT  -1.765000  32.655000  -1.595000  32.825000 ;
      RECT  -1.765000  33.875000  -1.595000  34.045000 ;
      RECT  -1.765000  35.095000  -1.595000  35.265000 ;
      RECT  -1.765000  36.315000  -1.595000  36.485000 ;
      RECT  -1.765000  37.535000  -1.595000  37.705000 ;
      RECT  -1.765000  38.755000  -1.595000  38.925000 ;
      RECT  -1.765000  39.975000  -1.595000  40.145000 ;
      RECT  -1.765000  41.195000  -1.595000  41.365000 ;
      RECT  -1.765000  42.415000  -1.595000  42.585000 ;
      RECT  -1.765000  43.635000  -1.595000  43.805000 ;
      RECT  -1.765000  44.855000  -1.595000  45.025000 ;
      RECT  -1.765000  46.075000  -1.595000  46.245000 ;
      RECT  -1.765000  47.295000  -1.595000  47.465000 ;
      RECT  -1.765000  48.515000  -1.595000  48.685000 ;
      RECT  -1.765000  49.735000  -1.595000  49.905000 ;
      RECT  -1.765000  50.955000  -1.595000  51.125000 ;
      RECT  -1.765000  52.175000  -1.595000  52.345000 ;
      RECT  -1.765000  53.395000  -1.595000  53.565000 ;
      RECT  -1.765000  54.615000  -1.595000  54.785000 ;
      RECT  -1.765000  55.835000  -1.595000  56.005000 ;
      RECT  -1.765000  57.055000  -1.595000  57.225000 ;
      RECT  -1.765000  58.275000  -1.595000  58.445000 ;
      RECT  -1.765000  59.495000  -1.595000  59.665000 ;
      RECT  -1.765000  60.715000  -1.595000  60.885000 ;
      RECT  -1.765000  61.935000  -1.595000  62.105000 ;
      RECT  -1.765000  63.155000  -1.595000  63.325000 ;
      RECT  -1.765000  64.375000  -1.595000  64.545000 ;
      RECT  -1.765000  65.595000  -1.595000  65.765000 ;
      RECT  -1.765000  66.815000  -1.595000  66.985000 ;
      RECT  -1.765000  68.035000  -1.595000  68.205000 ;
      RECT  -1.765000  69.255000  -1.595000  69.425000 ;
      RECT  -1.765000  70.475000  -1.595000  70.645000 ;
      RECT  -1.765000  71.695000  -1.595000  71.865000 ;
      RECT  -1.765000  72.915000  -1.595000  73.085000 ;
      RECT  -1.765000  74.135000  -1.595000  74.305000 ;
      RECT  -1.765000  75.355000  -1.595000  75.525000 ;
      RECT  -1.765000  76.575000  -1.595000  76.745000 ;
      RECT  -1.765000  77.795000  -1.595000  77.965000 ;
      RECT  -1.765000  79.015000  -1.595000  79.185000 ;
      RECT  -1.765000  80.235000  -1.595000  80.405000 ;
      RECT  -1.765000  81.455000  -1.595000  81.625000 ;
      RECT  -1.765000  82.675000  -1.595000  82.845000 ;
      RECT  -1.765000  83.895000  -1.595000  84.065000 ;
      RECT  -1.765000  85.115000  -1.595000  85.285000 ;
      RECT  -1.765000  86.335000  -1.595000  86.505000 ;
      RECT  -1.765000  87.555000  -1.595000  87.725000 ;
      RECT  -1.765000  88.775000  -1.595000  88.945000 ;
      RECT  -1.765000  89.995000  -1.595000  90.165000 ;
      RECT  -1.765000  91.215000  -1.595000  91.385000 ;
      RECT  -1.765000  92.435000  -1.595000  92.605000 ;
      RECT  -1.765000  93.655000  -1.595000  93.825000 ;
      RECT  -1.765000  94.875000  -1.595000  95.045000 ;
      RECT  -1.765000  96.095000  -1.595000  96.265000 ;
      RECT  -1.765000  97.315000  -1.595000  97.485000 ;
      RECT  -1.765000  98.535000  -1.595000  98.705000 ;
      RECT  -1.765000  99.755000  -1.595000  99.925000 ;
      RECT  -1.765000 100.975000  -1.595000 101.145000 ;
      RECT  -1.765000 102.195000  -1.595000 102.365000 ;
      RECT  -1.765000 103.415000  -1.595000 103.585000 ;
      RECT  -1.765000 104.635000  -1.595000 104.805000 ;
      RECT  -1.765000 105.855000  -1.595000 106.025000 ;
      RECT  -1.765000 107.075000  -1.595000 107.245000 ;
      RECT  -1.765000 108.295000  -1.595000 108.465000 ;
      RECT  -1.765000 109.515000  -1.595000 109.685000 ;
      RECT  -1.765000 110.735000  -1.595000 110.905000 ;
      RECT  -1.765000 111.955000  -1.595000 112.125000 ;
      RECT  -1.765000 113.175000  -1.595000 113.345000 ;
      RECT  -1.765000 114.395000  -1.595000 114.565000 ;
      RECT  -1.765000 115.615000  -1.595000 115.785000 ;
      RECT  -1.765000 116.835000  -1.595000 117.005000 ;
      RECT  -1.765000 118.055000  -1.595000 118.225000 ;
      RECT  -1.765000 119.275000  -1.595000 119.445000 ;
      RECT  -1.765000 120.495000  -1.595000 120.665000 ;
      RECT  -1.765000 121.715000  -1.595000 121.885000 ;
      RECT  -1.765000 122.935000  -1.595000 123.105000 ;
      RECT  -1.765000 124.155000  -1.595000 124.325000 ;
      RECT  -1.765000 125.375000  -1.595000 125.545000 ;
      RECT  -1.765000 126.595000  -1.595000 126.765000 ;
      RECT  -1.765000 127.815000  -1.595000 127.985000 ;
      RECT  -1.765000 129.035000  -1.595000 129.205000 ;
      RECT  -1.765000 130.255000  -1.595000 130.425000 ;
      RECT  -1.765000 131.475000  -1.595000 131.645000 ;
      RECT  -1.765000 132.695000  -1.595000 132.865000 ;
      RECT  -1.765000 133.915000  -1.595000 134.085000 ;
      RECT  -1.765000 135.135000  -1.595000 135.305000 ;
      RECT  -1.765000 136.355000  -1.595000 136.525000 ;
      RECT  -1.765000 137.575000  -1.595000 137.745000 ;
      RECT  -1.765000 138.795000  -1.595000 138.965000 ;
      RECT  -1.765000 140.015000  -1.595000 140.185000 ;
      RECT  -1.765000 141.235000  -1.595000 141.405000 ;
      RECT  -1.765000 142.455000  -1.595000 142.625000 ;
      RECT  -1.765000 143.675000  -1.595000 143.845000 ;
      RECT  -1.765000 144.895000  -1.595000 145.065000 ;
      RECT  -1.765000 146.115000  -1.595000 146.285000 ;
      RECT  -1.765000 147.335000  -1.595000 147.505000 ;
      RECT  -1.765000 148.555000  -1.595000 148.725000 ;
      RECT  -1.765000 149.775000  -1.595000 149.945000 ;
      RECT  -1.765000 150.995000  -1.595000 151.165000 ;
      RECT  -1.765000 152.215000  -1.595000 152.385000 ;
      RECT  -1.765000 153.435000  -1.595000 153.605000 ;
      RECT  -1.765000 154.655000  -1.595000 154.825000 ;
      RECT  -1.670000 156.415000  -1.500000 156.585000 ;
      RECT  -1.440000  -8.145000  -1.270000  -7.975000 ;
      RECT  -1.310000 156.415000  -1.140000 156.585000 ;
      RECT  -1.285000  -6.385000  -1.115000  -6.215000 ;
      RECT  -1.285000  -5.165000  -1.115000  -4.995000 ;
      RECT  -1.285000  -3.945000  -1.115000  -3.775000 ;
      RECT  -1.285000  -2.725000  -1.115000  -2.555000 ;
      RECT  -1.285000  -1.505000  -1.115000  -1.335000 ;
      RECT  -1.285000  -0.285000  -1.115000  -0.115000 ;
      RECT  -1.285000   0.935000  -1.115000   1.105000 ;
      RECT  -1.285000   2.155000  -1.115000   2.325000 ;
      RECT  -1.285000   3.375000  -1.115000   3.545000 ;
      RECT  -1.285000   4.595000  -1.115000   4.765000 ;
      RECT  -1.285000   5.815000  -1.115000   5.985000 ;
      RECT  -1.285000   7.035000  -1.115000   7.205000 ;
      RECT  -1.285000   8.255000  -1.115000   8.425000 ;
      RECT  -1.285000   9.475000  -1.115000   9.645000 ;
      RECT  -1.285000  10.695000  -1.115000  10.865000 ;
      RECT  -1.285000  11.915000  -1.115000  12.085000 ;
      RECT  -1.285000  13.135000  -1.115000  13.305000 ;
      RECT  -1.285000  14.355000  -1.115000  14.525000 ;
      RECT  -1.285000  15.575000  -1.115000  15.745000 ;
      RECT  -1.285000  16.795000  -1.115000  16.965000 ;
      RECT  -1.285000  18.015000  -1.115000  18.185000 ;
      RECT  -1.285000  19.235000  -1.115000  19.405000 ;
      RECT  -1.285000  20.455000  -1.115000  20.625000 ;
      RECT  -1.285000  21.675000  -1.115000  21.845000 ;
      RECT  -1.285000  22.895000  -1.115000  23.065000 ;
      RECT  -1.285000  24.115000  -1.115000  24.285000 ;
      RECT  -1.285000  25.335000  -1.115000  25.505000 ;
      RECT  -1.285000  26.555000  -1.115000  26.725000 ;
      RECT  -1.285000  27.775000  -1.115000  27.945000 ;
      RECT  -1.285000  28.995000  -1.115000  29.165000 ;
      RECT  -1.285000  30.215000  -1.115000  30.385000 ;
      RECT  -1.285000  31.435000  -1.115000  31.605000 ;
      RECT  -1.285000  32.655000  -1.115000  32.825000 ;
      RECT  -1.285000  33.875000  -1.115000  34.045000 ;
      RECT  -1.285000  35.095000  -1.115000  35.265000 ;
      RECT  -1.285000  36.315000  -1.115000  36.485000 ;
      RECT  -1.285000  37.535000  -1.115000  37.705000 ;
      RECT  -1.285000  38.755000  -1.115000  38.925000 ;
      RECT  -1.285000  39.975000  -1.115000  40.145000 ;
      RECT  -1.285000  41.195000  -1.115000  41.365000 ;
      RECT  -1.285000  42.415000  -1.115000  42.585000 ;
      RECT  -1.285000  43.635000  -1.115000  43.805000 ;
      RECT  -1.285000  44.855000  -1.115000  45.025000 ;
      RECT  -1.285000  46.075000  -1.115000  46.245000 ;
      RECT  -1.285000  47.295000  -1.115000  47.465000 ;
      RECT  -1.285000  48.515000  -1.115000  48.685000 ;
      RECT  -1.285000  49.735000  -1.115000  49.905000 ;
      RECT  -1.285000  50.955000  -1.115000  51.125000 ;
      RECT  -1.285000  52.175000  -1.115000  52.345000 ;
      RECT  -1.285000  53.395000  -1.115000  53.565000 ;
      RECT  -1.285000  54.615000  -1.115000  54.785000 ;
      RECT  -1.285000  55.835000  -1.115000  56.005000 ;
      RECT  -1.285000  57.055000  -1.115000  57.225000 ;
      RECT  -1.285000  58.275000  -1.115000  58.445000 ;
      RECT  -1.285000  59.495000  -1.115000  59.665000 ;
      RECT  -1.285000  60.715000  -1.115000  60.885000 ;
      RECT  -1.285000  61.935000  -1.115000  62.105000 ;
      RECT  -1.285000  63.155000  -1.115000  63.325000 ;
      RECT  -1.285000  64.375000  -1.115000  64.545000 ;
      RECT  -1.285000  65.595000  -1.115000  65.765000 ;
      RECT  -1.285000  66.815000  -1.115000  66.985000 ;
      RECT  -1.285000  68.035000  -1.115000  68.205000 ;
      RECT  -1.285000  69.255000  -1.115000  69.425000 ;
      RECT  -1.285000  70.475000  -1.115000  70.645000 ;
      RECT  -1.285000  71.695000  -1.115000  71.865000 ;
      RECT  -1.285000  72.915000  -1.115000  73.085000 ;
      RECT  -1.285000  74.135000  -1.115000  74.305000 ;
      RECT  -1.285000  75.355000  -1.115000  75.525000 ;
      RECT  -1.285000  76.575000  -1.115000  76.745000 ;
      RECT  -1.285000  77.795000  -1.115000  77.965000 ;
      RECT  -1.285000  79.015000  -1.115000  79.185000 ;
      RECT  -1.285000  80.235000  -1.115000  80.405000 ;
      RECT  -1.285000  81.455000  -1.115000  81.625000 ;
      RECT  -1.285000  82.675000  -1.115000  82.845000 ;
      RECT  -1.285000  83.895000  -1.115000  84.065000 ;
      RECT  -1.285000  85.115000  -1.115000  85.285000 ;
      RECT  -1.285000  86.335000  -1.115000  86.505000 ;
      RECT  -1.285000  87.555000  -1.115000  87.725000 ;
      RECT  -1.285000  88.775000  -1.115000  88.945000 ;
      RECT  -1.285000  89.995000  -1.115000  90.165000 ;
      RECT  -1.285000  91.215000  -1.115000  91.385000 ;
      RECT  -1.285000  92.435000  -1.115000  92.605000 ;
      RECT  -1.285000  93.655000  -1.115000  93.825000 ;
      RECT  -1.285000  94.875000  -1.115000  95.045000 ;
      RECT  -1.285000  96.095000  -1.115000  96.265000 ;
      RECT  -1.285000  97.315000  -1.115000  97.485000 ;
      RECT  -1.285000  98.535000  -1.115000  98.705000 ;
      RECT  -1.285000  99.755000  -1.115000  99.925000 ;
      RECT  -1.285000 100.975000  -1.115000 101.145000 ;
      RECT  -1.285000 102.195000  -1.115000 102.365000 ;
      RECT  -1.285000 103.415000  -1.115000 103.585000 ;
      RECT  -1.285000 104.635000  -1.115000 104.805000 ;
      RECT  -1.285000 105.855000  -1.115000 106.025000 ;
      RECT  -1.285000 107.075000  -1.115000 107.245000 ;
      RECT  -1.285000 108.295000  -1.115000 108.465000 ;
      RECT  -1.285000 109.515000  -1.115000 109.685000 ;
      RECT  -1.285000 110.735000  -1.115000 110.905000 ;
      RECT  -1.285000 111.955000  -1.115000 112.125000 ;
      RECT  -1.285000 113.175000  -1.115000 113.345000 ;
      RECT  -1.285000 114.395000  -1.115000 114.565000 ;
      RECT  -1.285000 115.615000  -1.115000 115.785000 ;
      RECT  -1.285000 116.835000  -1.115000 117.005000 ;
      RECT  -1.285000 118.055000  -1.115000 118.225000 ;
      RECT  -1.285000 119.275000  -1.115000 119.445000 ;
      RECT  -1.285000 120.495000  -1.115000 120.665000 ;
      RECT  -1.285000 121.715000  -1.115000 121.885000 ;
      RECT  -1.285000 122.935000  -1.115000 123.105000 ;
      RECT  -1.285000 124.155000  -1.115000 124.325000 ;
      RECT  -1.285000 125.375000  -1.115000 125.545000 ;
      RECT  -1.285000 126.595000  -1.115000 126.765000 ;
      RECT  -1.285000 127.815000  -1.115000 127.985000 ;
      RECT  -1.285000 129.035000  -1.115000 129.205000 ;
      RECT  -1.285000 130.255000  -1.115000 130.425000 ;
      RECT  -1.285000 131.475000  -1.115000 131.645000 ;
      RECT  -1.285000 132.695000  -1.115000 132.865000 ;
      RECT  -1.285000 133.915000  -1.115000 134.085000 ;
      RECT  -1.285000 135.135000  -1.115000 135.305000 ;
      RECT  -1.285000 136.355000  -1.115000 136.525000 ;
      RECT  -1.285000 137.575000  -1.115000 137.745000 ;
      RECT  -1.285000 138.795000  -1.115000 138.965000 ;
      RECT  -1.285000 140.015000  -1.115000 140.185000 ;
      RECT  -1.285000 141.235000  -1.115000 141.405000 ;
      RECT  -1.285000 142.455000  -1.115000 142.625000 ;
      RECT  -1.285000 143.675000  -1.115000 143.845000 ;
      RECT  -1.285000 144.895000  -1.115000 145.065000 ;
      RECT  -1.285000 146.115000  -1.115000 146.285000 ;
      RECT  -1.285000 147.335000  -1.115000 147.505000 ;
      RECT  -1.285000 148.555000  -1.115000 148.725000 ;
      RECT  -1.285000 149.775000  -1.115000 149.945000 ;
      RECT  -1.285000 150.995000  -1.115000 151.165000 ;
      RECT  -1.285000 152.215000  -1.115000 152.385000 ;
      RECT  -1.285000 153.435000  -1.115000 153.605000 ;
      RECT  -1.285000 154.655000  -1.115000 154.825000 ;
      RECT  -1.080000  -8.145000  -0.910000  -7.975000 ;
      RECT  -0.950000 156.415000  -0.780000 156.585000 ;
      RECT  -0.805000  -6.385000  -0.635000  -6.215000 ;
      RECT  -0.805000  -5.165000  -0.635000  -4.995000 ;
      RECT  -0.805000  -3.945000  -0.635000  -3.775000 ;
      RECT  -0.805000  -2.725000  -0.635000  -2.555000 ;
      RECT  -0.805000  -1.505000  -0.635000  -1.335000 ;
      RECT  -0.805000  -0.285000  -0.635000  -0.115000 ;
      RECT  -0.805000   0.935000  -0.635000   1.105000 ;
      RECT  -0.805000   2.155000  -0.635000   2.325000 ;
      RECT  -0.805000   3.375000  -0.635000   3.545000 ;
      RECT  -0.805000   4.595000  -0.635000   4.765000 ;
      RECT  -0.805000   5.815000  -0.635000   5.985000 ;
      RECT  -0.805000   7.035000  -0.635000   7.205000 ;
      RECT  -0.805000   8.255000  -0.635000   8.425000 ;
      RECT  -0.805000   9.475000  -0.635000   9.645000 ;
      RECT  -0.805000  10.695000  -0.635000  10.865000 ;
      RECT  -0.805000  11.915000  -0.635000  12.085000 ;
      RECT  -0.805000  13.135000  -0.635000  13.305000 ;
      RECT  -0.805000  14.355000  -0.635000  14.525000 ;
      RECT  -0.805000  15.575000  -0.635000  15.745000 ;
      RECT  -0.805000  16.795000  -0.635000  16.965000 ;
      RECT  -0.805000  18.015000  -0.635000  18.185000 ;
      RECT  -0.805000  19.235000  -0.635000  19.405000 ;
      RECT  -0.805000  20.455000  -0.635000  20.625000 ;
      RECT  -0.805000  21.675000  -0.635000  21.845000 ;
      RECT  -0.805000  22.895000  -0.635000  23.065000 ;
      RECT  -0.805000  24.115000  -0.635000  24.285000 ;
      RECT  -0.805000  25.335000  -0.635000  25.505000 ;
      RECT  -0.805000  26.555000  -0.635000  26.725000 ;
      RECT  -0.805000  27.775000  -0.635000  27.945000 ;
      RECT  -0.805000  28.995000  -0.635000  29.165000 ;
      RECT  -0.805000  30.215000  -0.635000  30.385000 ;
      RECT  -0.805000  31.435000  -0.635000  31.605000 ;
      RECT  -0.805000  32.655000  -0.635000  32.825000 ;
      RECT  -0.805000  33.875000  -0.635000  34.045000 ;
      RECT  -0.805000  35.095000  -0.635000  35.265000 ;
      RECT  -0.805000  36.315000  -0.635000  36.485000 ;
      RECT  -0.805000  37.535000  -0.635000  37.705000 ;
      RECT  -0.805000  38.755000  -0.635000  38.925000 ;
      RECT  -0.805000  39.975000  -0.635000  40.145000 ;
      RECT  -0.805000  41.195000  -0.635000  41.365000 ;
      RECT  -0.805000  42.415000  -0.635000  42.585000 ;
      RECT  -0.805000  43.635000  -0.635000  43.805000 ;
      RECT  -0.805000  44.855000  -0.635000  45.025000 ;
      RECT  -0.805000  46.075000  -0.635000  46.245000 ;
      RECT  -0.805000  47.295000  -0.635000  47.465000 ;
      RECT  -0.805000  48.515000  -0.635000  48.685000 ;
      RECT  -0.805000  49.735000  -0.635000  49.905000 ;
      RECT  -0.805000  50.955000  -0.635000  51.125000 ;
      RECT  -0.805000  52.175000  -0.635000  52.345000 ;
      RECT  -0.805000  53.395000  -0.635000  53.565000 ;
      RECT  -0.805000  54.615000  -0.635000  54.785000 ;
      RECT  -0.805000  55.835000  -0.635000  56.005000 ;
      RECT  -0.805000  57.055000  -0.635000  57.225000 ;
      RECT  -0.805000  58.275000  -0.635000  58.445000 ;
      RECT  -0.805000  59.495000  -0.635000  59.665000 ;
      RECT  -0.805000  60.715000  -0.635000  60.885000 ;
      RECT  -0.805000  61.935000  -0.635000  62.105000 ;
      RECT  -0.805000  63.155000  -0.635000  63.325000 ;
      RECT  -0.805000  64.375000  -0.635000  64.545000 ;
      RECT  -0.805000  65.595000  -0.635000  65.765000 ;
      RECT  -0.805000  66.815000  -0.635000  66.985000 ;
      RECT  -0.805000  68.035000  -0.635000  68.205000 ;
      RECT  -0.805000  69.255000  -0.635000  69.425000 ;
      RECT  -0.805000  70.475000  -0.635000  70.645000 ;
      RECT  -0.805000  71.695000  -0.635000  71.865000 ;
      RECT  -0.805000  72.915000  -0.635000  73.085000 ;
      RECT  -0.805000  74.135000  -0.635000  74.305000 ;
      RECT  -0.805000  75.355000  -0.635000  75.525000 ;
      RECT  -0.805000  76.575000  -0.635000  76.745000 ;
      RECT  -0.805000  77.795000  -0.635000  77.965000 ;
      RECT  -0.805000  79.015000  -0.635000  79.185000 ;
      RECT  -0.805000  80.235000  -0.635000  80.405000 ;
      RECT  -0.805000  81.455000  -0.635000  81.625000 ;
      RECT  -0.805000  82.675000  -0.635000  82.845000 ;
      RECT  -0.805000  83.895000  -0.635000  84.065000 ;
      RECT  -0.805000  85.115000  -0.635000  85.285000 ;
      RECT  -0.805000  86.335000  -0.635000  86.505000 ;
      RECT  -0.805000  87.555000  -0.635000  87.725000 ;
      RECT  -0.805000  88.775000  -0.635000  88.945000 ;
      RECT  -0.805000  89.995000  -0.635000  90.165000 ;
      RECT  -0.805000  91.215000  -0.635000  91.385000 ;
      RECT  -0.805000  92.435000  -0.635000  92.605000 ;
      RECT  -0.805000  93.655000  -0.635000  93.825000 ;
      RECT  -0.805000  94.875000  -0.635000  95.045000 ;
      RECT  -0.805000  96.095000  -0.635000  96.265000 ;
      RECT  -0.805000  97.315000  -0.635000  97.485000 ;
      RECT  -0.805000  98.535000  -0.635000  98.705000 ;
      RECT  -0.805000  99.755000  -0.635000  99.925000 ;
      RECT  -0.805000 100.975000  -0.635000 101.145000 ;
      RECT  -0.805000 102.195000  -0.635000 102.365000 ;
      RECT  -0.805000 103.415000  -0.635000 103.585000 ;
      RECT  -0.805000 104.635000  -0.635000 104.805000 ;
      RECT  -0.805000 105.855000  -0.635000 106.025000 ;
      RECT  -0.805000 107.075000  -0.635000 107.245000 ;
      RECT  -0.805000 108.295000  -0.635000 108.465000 ;
      RECT  -0.805000 109.515000  -0.635000 109.685000 ;
      RECT  -0.805000 110.735000  -0.635000 110.905000 ;
      RECT  -0.805000 111.955000  -0.635000 112.125000 ;
      RECT  -0.805000 113.175000  -0.635000 113.345000 ;
      RECT  -0.805000 114.395000  -0.635000 114.565000 ;
      RECT  -0.805000 115.615000  -0.635000 115.785000 ;
      RECT  -0.805000 116.835000  -0.635000 117.005000 ;
      RECT  -0.805000 118.055000  -0.635000 118.225000 ;
      RECT  -0.805000 119.275000  -0.635000 119.445000 ;
      RECT  -0.805000 120.495000  -0.635000 120.665000 ;
      RECT  -0.805000 121.715000  -0.635000 121.885000 ;
      RECT  -0.805000 122.935000  -0.635000 123.105000 ;
      RECT  -0.805000 124.155000  -0.635000 124.325000 ;
      RECT  -0.805000 125.375000  -0.635000 125.545000 ;
      RECT  -0.805000 126.595000  -0.635000 126.765000 ;
      RECT  -0.805000 127.815000  -0.635000 127.985000 ;
      RECT  -0.805000 129.035000  -0.635000 129.205000 ;
      RECT  -0.805000 130.255000  -0.635000 130.425000 ;
      RECT  -0.805000 131.475000  -0.635000 131.645000 ;
      RECT  -0.805000 132.695000  -0.635000 132.865000 ;
      RECT  -0.805000 133.915000  -0.635000 134.085000 ;
      RECT  -0.805000 135.135000  -0.635000 135.305000 ;
      RECT  -0.805000 136.355000  -0.635000 136.525000 ;
      RECT  -0.805000 137.575000  -0.635000 137.745000 ;
      RECT  -0.805000 138.795000  -0.635000 138.965000 ;
      RECT  -0.805000 140.015000  -0.635000 140.185000 ;
      RECT  -0.805000 141.235000  -0.635000 141.405000 ;
      RECT  -0.805000 142.455000  -0.635000 142.625000 ;
      RECT  -0.805000 143.675000  -0.635000 143.845000 ;
      RECT  -0.805000 144.895000  -0.635000 145.065000 ;
      RECT  -0.805000 146.115000  -0.635000 146.285000 ;
      RECT  -0.805000 147.335000  -0.635000 147.505000 ;
      RECT  -0.805000 148.555000  -0.635000 148.725000 ;
      RECT  -0.805000 149.775000  -0.635000 149.945000 ;
      RECT  -0.805000 150.995000  -0.635000 151.165000 ;
      RECT  -0.805000 152.215000  -0.635000 152.385000 ;
      RECT  -0.805000 153.435000  -0.635000 153.605000 ;
      RECT  -0.805000 154.655000  -0.635000 154.825000 ;
      RECT  -0.720000  -8.145000  -0.550000  -7.975000 ;
      RECT  -0.590000 156.415000  -0.420000 156.585000 ;
      RECT  -0.360000  -8.145000  -0.190000  -7.975000 ;
      RECT  -0.325000  -6.385000  -0.155000  -6.215000 ;
      RECT  -0.325000  -5.165000  -0.155000  -4.995000 ;
      RECT  -0.325000  -3.945000  -0.155000  -3.775000 ;
      RECT  -0.325000  -2.725000  -0.155000  -2.555000 ;
      RECT  -0.325000  -1.505000  -0.155000  -1.335000 ;
      RECT  -0.325000  -0.285000  -0.155000  -0.115000 ;
      RECT  -0.325000   0.935000  -0.155000   1.105000 ;
      RECT  -0.325000   2.155000  -0.155000   2.325000 ;
      RECT  -0.325000   3.375000  -0.155000   3.545000 ;
      RECT  -0.325000   4.595000  -0.155000   4.765000 ;
      RECT  -0.325000   5.815000  -0.155000   5.985000 ;
      RECT  -0.325000   7.035000  -0.155000   7.205000 ;
      RECT  -0.325000   8.255000  -0.155000   8.425000 ;
      RECT  -0.325000   9.475000  -0.155000   9.645000 ;
      RECT  -0.325000  10.695000  -0.155000  10.865000 ;
      RECT  -0.325000  11.915000  -0.155000  12.085000 ;
      RECT  -0.325000  13.135000  -0.155000  13.305000 ;
      RECT  -0.325000  14.355000  -0.155000  14.525000 ;
      RECT  -0.325000  15.575000  -0.155000  15.745000 ;
      RECT  -0.325000  16.795000  -0.155000  16.965000 ;
      RECT  -0.325000  18.015000  -0.155000  18.185000 ;
      RECT  -0.325000  19.235000  -0.155000  19.405000 ;
      RECT  -0.325000  20.455000  -0.155000  20.625000 ;
      RECT  -0.325000  21.675000  -0.155000  21.845000 ;
      RECT  -0.325000  22.895000  -0.155000  23.065000 ;
      RECT  -0.325000  24.115000  -0.155000  24.285000 ;
      RECT  -0.325000  25.335000  -0.155000  25.505000 ;
      RECT  -0.325000  26.555000  -0.155000  26.725000 ;
      RECT  -0.325000  27.775000  -0.155000  27.945000 ;
      RECT  -0.325000  28.995000  -0.155000  29.165000 ;
      RECT  -0.325000  30.215000  -0.155000  30.385000 ;
      RECT  -0.325000  31.435000  -0.155000  31.605000 ;
      RECT  -0.325000  32.655000  -0.155000  32.825000 ;
      RECT  -0.325000  33.875000  -0.155000  34.045000 ;
      RECT  -0.325000  35.095000  -0.155000  35.265000 ;
      RECT  -0.325000  36.315000  -0.155000  36.485000 ;
      RECT  -0.325000  37.535000  -0.155000  37.705000 ;
      RECT  -0.325000  38.755000  -0.155000  38.925000 ;
      RECT  -0.325000  39.975000  -0.155000  40.145000 ;
      RECT  -0.325000  41.195000  -0.155000  41.365000 ;
      RECT  -0.325000  42.415000  -0.155000  42.585000 ;
      RECT  -0.325000  43.635000  -0.155000  43.805000 ;
      RECT  -0.325000  44.855000  -0.155000  45.025000 ;
      RECT  -0.325000  46.075000  -0.155000  46.245000 ;
      RECT  -0.325000  47.295000  -0.155000  47.465000 ;
      RECT  -0.325000  48.515000  -0.155000  48.685000 ;
      RECT  -0.325000  49.735000  -0.155000  49.905000 ;
      RECT  -0.325000  50.955000  -0.155000  51.125000 ;
      RECT  -0.325000  52.175000  -0.155000  52.345000 ;
      RECT  -0.325000  53.395000  -0.155000  53.565000 ;
      RECT  -0.325000  54.615000  -0.155000  54.785000 ;
      RECT  -0.325000  55.835000  -0.155000  56.005000 ;
      RECT  -0.325000  57.055000  -0.155000  57.225000 ;
      RECT  -0.325000  58.275000  -0.155000  58.445000 ;
      RECT  -0.325000  59.495000  -0.155000  59.665000 ;
      RECT  -0.325000  60.715000  -0.155000  60.885000 ;
      RECT  -0.325000  61.935000  -0.155000  62.105000 ;
      RECT  -0.325000  63.155000  -0.155000  63.325000 ;
      RECT  -0.325000  64.375000  -0.155000  64.545000 ;
      RECT  -0.325000  65.595000  -0.155000  65.765000 ;
      RECT  -0.325000  66.815000  -0.155000  66.985000 ;
      RECT  -0.325000  68.035000  -0.155000  68.205000 ;
      RECT  -0.325000  69.255000  -0.155000  69.425000 ;
      RECT  -0.325000  70.475000  -0.155000  70.645000 ;
      RECT  -0.325000  71.695000  -0.155000  71.865000 ;
      RECT  -0.325000  72.915000  -0.155000  73.085000 ;
      RECT  -0.325000  74.135000  -0.155000  74.305000 ;
      RECT  -0.325000  75.355000  -0.155000  75.525000 ;
      RECT  -0.325000  76.575000  -0.155000  76.745000 ;
      RECT  -0.325000  77.795000  -0.155000  77.965000 ;
      RECT  -0.325000  79.015000  -0.155000  79.185000 ;
      RECT  -0.325000  80.235000  -0.155000  80.405000 ;
      RECT  -0.325000  81.455000  -0.155000  81.625000 ;
      RECT  -0.325000  82.675000  -0.155000  82.845000 ;
      RECT  -0.325000  83.895000  -0.155000  84.065000 ;
      RECT  -0.325000  85.115000  -0.155000  85.285000 ;
      RECT  -0.325000  86.335000  -0.155000  86.505000 ;
      RECT  -0.325000  87.555000  -0.155000  87.725000 ;
      RECT  -0.325000  88.775000  -0.155000  88.945000 ;
      RECT  -0.325000  89.995000  -0.155000  90.165000 ;
      RECT  -0.325000  91.215000  -0.155000  91.385000 ;
      RECT  -0.325000  92.435000  -0.155000  92.605000 ;
      RECT  -0.325000  93.655000  -0.155000  93.825000 ;
      RECT  -0.325000  94.875000  -0.155000  95.045000 ;
      RECT  -0.325000  96.095000  -0.155000  96.265000 ;
      RECT  -0.325000  97.315000  -0.155000  97.485000 ;
      RECT  -0.325000  98.535000  -0.155000  98.705000 ;
      RECT  -0.325000  99.755000  -0.155000  99.925000 ;
      RECT  -0.325000 100.975000  -0.155000 101.145000 ;
      RECT  -0.325000 102.195000  -0.155000 102.365000 ;
      RECT  -0.325000 103.415000  -0.155000 103.585000 ;
      RECT  -0.325000 104.635000  -0.155000 104.805000 ;
      RECT  -0.325000 105.855000  -0.155000 106.025000 ;
      RECT  -0.325000 107.075000  -0.155000 107.245000 ;
      RECT  -0.325000 108.295000  -0.155000 108.465000 ;
      RECT  -0.325000 109.515000  -0.155000 109.685000 ;
      RECT  -0.325000 110.735000  -0.155000 110.905000 ;
      RECT  -0.325000 111.955000  -0.155000 112.125000 ;
      RECT  -0.325000 113.175000  -0.155000 113.345000 ;
      RECT  -0.325000 114.395000  -0.155000 114.565000 ;
      RECT  -0.325000 115.615000  -0.155000 115.785000 ;
      RECT  -0.325000 116.835000  -0.155000 117.005000 ;
      RECT  -0.325000 118.055000  -0.155000 118.225000 ;
      RECT  -0.325000 119.275000  -0.155000 119.445000 ;
      RECT  -0.325000 120.495000  -0.155000 120.665000 ;
      RECT  -0.325000 121.715000  -0.155000 121.885000 ;
      RECT  -0.325000 122.935000  -0.155000 123.105000 ;
      RECT  -0.325000 124.155000  -0.155000 124.325000 ;
      RECT  -0.325000 125.375000  -0.155000 125.545000 ;
      RECT  -0.325000 126.595000  -0.155000 126.765000 ;
      RECT  -0.325000 127.815000  -0.155000 127.985000 ;
      RECT  -0.325000 129.035000  -0.155000 129.205000 ;
      RECT  -0.325000 130.255000  -0.155000 130.425000 ;
      RECT  -0.325000 131.475000  -0.155000 131.645000 ;
      RECT  -0.325000 132.695000  -0.155000 132.865000 ;
      RECT  -0.325000 133.915000  -0.155000 134.085000 ;
      RECT  -0.325000 135.135000  -0.155000 135.305000 ;
      RECT  -0.325000 136.355000  -0.155000 136.525000 ;
      RECT  -0.325000 137.575000  -0.155000 137.745000 ;
      RECT  -0.325000 138.795000  -0.155000 138.965000 ;
      RECT  -0.325000 140.015000  -0.155000 140.185000 ;
      RECT  -0.325000 141.235000  -0.155000 141.405000 ;
      RECT  -0.325000 142.455000  -0.155000 142.625000 ;
      RECT  -0.325000 143.675000  -0.155000 143.845000 ;
      RECT  -0.325000 144.895000  -0.155000 145.065000 ;
      RECT  -0.325000 146.115000  -0.155000 146.285000 ;
      RECT  -0.325000 147.335000  -0.155000 147.505000 ;
      RECT  -0.325000 148.555000  -0.155000 148.725000 ;
      RECT  -0.325000 149.775000  -0.155000 149.945000 ;
      RECT  -0.325000 150.995000  -0.155000 151.165000 ;
      RECT  -0.325000 152.215000  -0.155000 152.385000 ;
      RECT  -0.325000 153.435000  -0.155000 153.605000 ;
      RECT  -0.325000 154.655000  -0.155000 154.825000 ;
      RECT  -0.230000 156.415000  -0.060000 156.585000 ;
      RECT   0.130000 156.415000   0.300000 156.585000 ;
      RECT   0.155000  -6.385000   0.325000  -6.215000 ;
      RECT   0.155000  -5.165000   0.325000  -4.995000 ;
      RECT   0.155000  -3.945000   0.325000  -3.775000 ;
      RECT   0.155000  -2.725000   0.325000  -2.555000 ;
      RECT   0.155000  -1.505000   0.325000  -1.335000 ;
      RECT   0.155000  -0.285000   0.325000  -0.115000 ;
      RECT   0.155000   0.935000   0.325000   1.105000 ;
      RECT   0.155000   2.155000   0.325000   2.325000 ;
      RECT   0.155000   3.375000   0.325000   3.545000 ;
      RECT   0.155000   4.595000   0.325000   4.765000 ;
      RECT   0.155000   5.815000   0.325000   5.985000 ;
      RECT   0.155000   7.035000   0.325000   7.205000 ;
      RECT   0.155000   8.255000   0.325000   8.425000 ;
      RECT   0.155000   9.475000   0.325000   9.645000 ;
      RECT   0.155000  10.695000   0.325000  10.865000 ;
      RECT   0.155000  11.915000   0.325000  12.085000 ;
      RECT   0.155000  13.135000   0.325000  13.305000 ;
      RECT   0.155000  14.355000   0.325000  14.525000 ;
      RECT   0.155000  15.575000   0.325000  15.745000 ;
      RECT   0.155000  16.795000   0.325000  16.965000 ;
      RECT   0.155000  18.015000   0.325000  18.185000 ;
      RECT   0.155000  19.235000   0.325000  19.405000 ;
      RECT   0.155000  20.455000   0.325000  20.625000 ;
      RECT   0.155000  21.675000   0.325000  21.845000 ;
      RECT   0.155000  22.895000   0.325000  23.065000 ;
      RECT   0.155000  24.115000   0.325000  24.285000 ;
      RECT   0.155000  25.335000   0.325000  25.505000 ;
      RECT   0.155000  26.555000   0.325000  26.725000 ;
      RECT   0.155000  27.775000   0.325000  27.945000 ;
      RECT   0.155000  28.995000   0.325000  29.165000 ;
      RECT   0.155000  30.215000   0.325000  30.385000 ;
      RECT   0.155000  31.435000   0.325000  31.605000 ;
      RECT   0.155000  32.655000   0.325000  32.825000 ;
      RECT   0.155000  33.875000   0.325000  34.045000 ;
      RECT   0.155000  35.095000   0.325000  35.265000 ;
      RECT   0.155000  36.315000   0.325000  36.485000 ;
      RECT   0.155000  37.535000   0.325000  37.705000 ;
      RECT   0.155000  38.755000   0.325000  38.925000 ;
      RECT   0.155000  39.975000   0.325000  40.145000 ;
      RECT   0.155000  41.195000   0.325000  41.365000 ;
      RECT   0.155000  42.415000   0.325000  42.585000 ;
      RECT   0.155000  43.635000   0.325000  43.805000 ;
      RECT   0.155000  44.855000   0.325000  45.025000 ;
      RECT   0.155000  46.075000   0.325000  46.245000 ;
      RECT   0.155000  47.295000   0.325000  47.465000 ;
      RECT   0.155000  48.515000   0.325000  48.685000 ;
      RECT   0.155000  49.735000   0.325000  49.905000 ;
      RECT   0.155000  50.955000   0.325000  51.125000 ;
      RECT   0.155000  52.175000   0.325000  52.345000 ;
      RECT   0.155000  53.395000   0.325000  53.565000 ;
      RECT   0.155000  54.615000   0.325000  54.785000 ;
      RECT   0.155000  55.835000   0.325000  56.005000 ;
      RECT   0.155000  57.055000   0.325000  57.225000 ;
      RECT   0.155000  58.275000   0.325000  58.445000 ;
      RECT   0.155000  59.495000   0.325000  59.665000 ;
      RECT   0.155000  60.715000   0.325000  60.885000 ;
      RECT   0.155000  61.935000   0.325000  62.105000 ;
      RECT   0.155000  63.155000   0.325000  63.325000 ;
      RECT   0.155000  64.375000   0.325000  64.545000 ;
      RECT   0.155000  65.595000   0.325000  65.765000 ;
      RECT   0.155000  66.815000   0.325000  66.985000 ;
      RECT   0.155000  68.035000   0.325000  68.205000 ;
      RECT   0.155000  69.255000   0.325000  69.425000 ;
      RECT   0.155000  70.475000   0.325000  70.645000 ;
      RECT   0.155000  71.695000   0.325000  71.865000 ;
      RECT   0.155000  72.915000   0.325000  73.085000 ;
      RECT   0.155000  74.135000   0.325000  74.305000 ;
      RECT   0.155000  75.355000   0.325000  75.525000 ;
      RECT   0.155000  76.575000   0.325000  76.745000 ;
      RECT   0.155000  77.795000   0.325000  77.965000 ;
      RECT   0.155000  79.015000   0.325000  79.185000 ;
      RECT   0.155000  80.235000   0.325000  80.405000 ;
      RECT   0.155000  81.455000   0.325000  81.625000 ;
      RECT   0.155000  82.675000   0.325000  82.845000 ;
      RECT   0.155000  83.895000   0.325000  84.065000 ;
      RECT   0.155000  85.115000   0.325000  85.285000 ;
      RECT   0.155000  86.335000   0.325000  86.505000 ;
      RECT   0.155000  87.555000   0.325000  87.725000 ;
      RECT   0.155000  88.775000   0.325000  88.945000 ;
      RECT   0.155000  89.995000   0.325000  90.165000 ;
      RECT   0.155000  91.215000   0.325000  91.385000 ;
      RECT   0.155000  92.435000   0.325000  92.605000 ;
      RECT   0.155000  93.655000   0.325000  93.825000 ;
      RECT   0.155000  94.875000   0.325000  95.045000 ;
      RECT   0.155000  96.095000   0.325000  96.265000 ;
      RECT   0.155000  97.315000   0.325000  97.485000 ;
      RECT   0.155000  98.535000   0.325000  98.705000 ;
      RECT   0.155000  99.755000   0.325000  99.925000 ;
      RECT   0.155000 100.975000   0.325000 101.145000 ;
      RECT   0.155000 102.195000   0.325000 102.365000 ;
      RECT   0.155000 103.415000   0.325000 103.585000 ;
      RECT   0.155000 104.635000   0.325000 104.805000 ;
      RECT   0.155000 105.855000   0.325000 106.025000 ;
      RECT   0.155000 107.075000   0.325000 107.245000 ;
      RECT   0.155000 108.295000   0.325000 108.465000 ;
      RECT   0.155000 109.515000   0.325000 109.685000 ;
      RECT   0.155000 110.735000   0.325000 110.905000 ;
      RECT   0.155000 111.955000   0.325000 112.125000 ;
      RECT   0.155000 113.175000   0.325000 113.345000 ;
      RECT   0.155000 114.395000   0.325000 114.565000 ;
      RECT   0.155000 115.615000   0.325000 115.785000 ;
      RECT   0.155000 116.835000   0.325000 117.005000 ;
      RECT   0.155000 118.055000   0.325000 118.225000 ;
      RECT   0.155000 119.275000   0.325000 119.445000 ;
      RECT   0.155000 120.495000   0.325000 120.665000 ;
      RECT   0.155000 121.715000   0.325000 121.885000 ;
      RECT   0.155000 122.935000   0.325000 123.105000 ;
      RECT   0.155000 124.155000   0.325000 124.325000 ;
      RECT   0.155000 125.375000   0.325000 125.545000 ;
      RECT   0.155000 126.595000   0.325000 126.765000 ;
      RECT   0.155000 127.815000   0.325000 127.985000 ;
      RECT   0.155000 129.035000   0.325000 129.205000 ;
      RECT   0.155000 130.255000   0.325000 130.425000 ;
      RECT   0.155000 131.475000   0.325000 131.645000 ;
      RECT   0.155000 132.695000   0.325000 132.865000 ;
      RECT   0.155000 133.915000   0.325000 134.085000 ;
      RECT   0.155000 135.135000   0.325000 135.305000 ;
      RECT   0.155000 136.355000   0.325000 136.525000 ;
      RECT   0.155000 137.575000   0.325000 137.745000 ;
      RECT   0.155000 138.795000   0.325000 138.965000 ;
      RECT   0.155000 140.015000   0.325000 140.185000 ;
      RECT   0.155000 141.235000   0.325000 141.405000 ;
      RECT   0.155000 142.455000   0.325000 142.625000 ;
      RECT   0.155000 143.675000   0.325000 143.845000 ;
      RECT   0.155000 144.895000   0.325000 145.065000 ;
      RECT   0.155000 146.115000   0.325000 146.285000 ;
      RECT   0.155000 147.335000   0.325000 147.505000 ;
      RECT   0.155000 148.555000   0.325000 148.725000 ;
      RECT   0.155000 149.775000   0.325000 149.945000 ;
      RECT   0.155000 150.995000   0.325000 151.165000 ;
      RECT   0.155000 152.215000   0.325000 152.385000 ;
      RECT   0.155000 153.435000   0.325000 153.605000 ;
      RECT   0.155000 154.655000   0.325000 154.825000 ;
      RECT   0.190000  -8.145000   0.360000  -7.975000 ;
      RECT   0.490000 156.415000   0.660000 156.585000 ;
      RECT   0.555000  -8.145000   0.725000  -7.975000 ;
      RECT   0.635000  -6.385000   0.805000  -6.215000 ;
      RECT   0.635000  -5.165000   0.805000  -4.995000 ;
      RECT   0.635000  -3.945000   0.805000  -3.775000 ;
      RECT   0.635000  -2.725000   0.805000  -2.555000 ;
      RECT   0.635000  -1.505000   0.805000  -1.335000 ;
      RECT   0.635000  -0.285000   0.805000  -0.115000 ;
      RECT   0.635000   0.935000   0.805000   1.105000 ;
      RECT   0.635000   2.155000   0.805000   2.325000 ;
      RECT   0.635000   3.375000   0.805000   3.545000 ;
      RECT   0.635000   4.595000   0.805000   4.765000 ;
      RECT   0.635000   5.815000   0.805000   5.985000 ;
      RECT   0.635000   7.035000   0.805000   7.205000 ;
      RECT   0.635000   8.255000   0.805000   8.425000 ;
      RECT   0.635000   9.475000   0.805000   9.645000 ;
      RECT   0.635000  10.695000   0.805000  10.865000 ;
      RECT   0.635000  11.915000   0.805000  12.085000 ;
      RECT   0.635000  13.135000   0.805000  13.305000 ;
      RECT   0.635000  14.355000   0.805000  14.525000 ;
      RECT   0.635000  15.575000   0.805000  15.745000 ;
      RECT   0.635000  16.795000   0.805000  16.965000 ;
      RECT   0.635000  18.015000   0.805000  18.185000 ;
      RECT   0.635000  19.235000   0.805000  19.405000 ;
      RECT   0.635000  20.455000   0.805000  20.625000 ;
      RECT   0.635000  21.675000   0.805000  21.845000 ;
      RECT   0.635000  22.895000   0.805000  23.065000 ;
      RECT   0.635000  24.115000   0.805000  24.285000 ;
      RECT   0.635000  25.335000   0.805000  25.505000 ;
      RECT   0.635000  26.555000   0.805000  26.725000 ;
      RECT   0.635000  27.775000   0.805000  27.945000 ;
      RECT   0.635000  28.995000   0.805000  29.165000 ;
      RECT   0.635000  30.215000   0.805000  30.385000 ;
      RECT   0.635000  31.435000   0.805000  31.605000 ;
      RECT   0.635000  32.655000   0.805000  32.825000 ;
      RECT   0.635000  33.875000   0.805000  34.045000 ;
      RECT   0.635000  35.095000   0.805000  35.265000 ;
      RECT   0.635000  36.315000   0.805000  36.485000 ;
      RECT   0.635000  37.535000   0.805000  37.705000 ;
      RECT   0.635000  38.755000   0.805000  38.925000 ;
      RECT   0.635000  39.975000   0.805000  40.145000 ;
      RECT   0.635000  41.195000   0.805000  41.365000 ;
      RECT   0.635000  42.415000   0.805000  42.585000 ;
      RECT   0.635000  43.635000   0.805000  43.805000 ;
      RECT   0.635000  44.855000   0.805000  45.025000 ;
      RECT   0.635000  46.075000   0.805000  46.245000 ;
      RECT   0.635000  47.295000   0.805000  47.465000 ;
      RECT   0.635000  48.515000   0.805000  48.685000 ;
      RECT   0.635000  49.735000   0.805000  49.905000 ;
      RECT   0.635000  50.955000   0.805000  51.125000 ;
      RECT   0.635000  52.175000   0.805000  52.345000 ;
      RECT   0.635000  53.395000   0.805000  53.565000 ;
      RECT   0.635000  54.615000   0.805000  54.785000 ;
      RECT   0.635000  55.835000   0.805000  56.005000 ;
      RECT   0.635000  57.055000   0.805000  57.225000 ;
      RECT   0.635000  58.275000   0.805000  58.445000 ;
      RECT   0.635000  59.495000   0.805000  59.665000 ;
      RECT   0.635000  60.715000   0.805000  60.885000 ;
      RECT   0.635000  61.935000   0.805000  62.105000 ;
      RECT   0.635000  63.155000   0.805000  63.325000 ;
      RECT   0.635000  64.375000   0.805000  64.545000 ;
      RECT   0.635000  65.595000   0.805000  65.765000 ;
      RECT   0.635000  66.815000   0.805000  66.985000 ;
      RECT   0.635000  68.035000   0.805000  68.205000 ;
      RECT   0.635000  69.255000   0.805000  69.425000 ;
      RECT   0.635000  70.475000   0.805000  70.645000 ;
      RECT   0.635000  71.695000   0.805000  71.865000 ;
      RECT   0.635000  72.915000   0.805000  73.085000 ;
      RECT   0.635000  74.135000   0.805000  74.305000 ;
      RECT   0.635000  75.355000   0.805000  75.525000 ;
      RECT   0.635000  76.575000   0.805000  76.745000 ;
      RECT   0.635000  77.795000   0.805000  77.965000 ;
      RECT   0.635000  79.015000   0.805000  79.185000 ;
      RECT   0.635000  80.235000   0.805000  80.405000 ;
      RECT   0.635000  81.455000   0.805000  81.625000 ;
      RECT   0.635000  82.675000   0.805000  82.845000 ;
      RECT   0.635000  83.895000   0.805000  84.065000 ;
      RECT   0.635000  85.115000   0.805000  85.285000 ;
      RECT   0.635000  86.335000   0.805000  86.505000 ;
      RECT   0.635000  87.555000   0.805000  87.725000 ;
      RECT   0.635000  88.775000   0.805000  88.945000 ;
      RECT   0.635000  89.995000   0.805000  90.165000 ;
      RECT   0.635000  91.215000   0.805000  91.385000 ;
      RECT   0.635000  92.435000   0.805000  92.605000 ;
      RECT   0.635000  93.655000   0.805000  93.825000 ;
      RECT   0.635000  94.875000   0.805000  95.045000 ;
      RECT   0.635000  96.095000   0.805000  96.265000 ;
      RECT   0.635000  97.315000   0.805000  97.485000 ;
      RECT   0.635000  98.535000   0.805000  98.705000 ;
      RECT   0.635000  99.755000   0.805000  99.925000 ;
      RECT   0.635000 100.975000   0.805000 101.145000 ;
      RECT   0.635000 102.195000   0.805000 102.365000 ;
      RECT   0.635000 103.415000   0.805000 103.585000 ;
      RECT   0.635000 104.635000   0.805000 104.805000 ;
      RECT   0.635000 105.855000   0.805000 106.025000 ;
      RECT   0.635000 107.075000   0.805000 107.245000 ;
      RECT   0.635000 108.295000   0.805000 108.465000 ;
      RECT   0.635000 109.515000   0.805000 109.685000 ;
      RECT   0.635000 110.735000   0.805000 110.905000 ;
      RECT   0.635000 111.955000   0.805000 112.125000 ;
      RECT   0.635000 113.175000   0.805000 113.345000 ;
      RECT   0.635000 114.395000   0.805000 114.565000 ;
      RECT   0.635000 115.615000   0.805000 115.785000 ;
      RECT   0.635000 116.835000   0.805000 117.005000 ;
      RECT   0.635000 118.055000   0.805000 118.225000 ;
      RECT   0.635000 119.275000   0.805000 119.445000 ;
      RECT   0.635000 120.495000   0.805000 120.665000 ;
      RECT   0.635000 121.715000   0.805000 121.885000 ;
      RECT   0.635000 122.935000   0.805000 123.105000 ;
      RECT   0.635000 124.155000   0.805000 124.325000 ;
      RECT   0.635000 125.375000   0.805000 125.545000 ;
      RECT   0.635000 126.595000   0.805000 126.765000 ;
      RECT   0.635000 127.815000   0.805000 127.985000 ;
      RECT   0.635000 129.035000   0.805000 129.205000 ;
      RECT   0.635000 130.255000   0.805000 130.425000 ;
      RECT   0.635000 131.475000   0.805000 131.645000 ;
      RECT   0.635000 132.695000   0.805000 132.865000 ;
      RECT   0.635000 133.915000   0.805000 134.085000 ;
      RECT   0.635000 135.135000   0.805000 135.305000 ;
      RECT   0.635000 136.355000   0.805000 136.525000 ;
      RECT   0.635000 137.575000   0.805000 137.745000 ;
      RECT   0.635000 138.795000   0.805000 138.965000 ;
      RECT   0.635000 140.015000   0.805000 140.185000 ;
      RECT   0.635000 141.235000   0.805000 141.405000 ;
      RECT   0.635000 142.455000   0.805000 142.625000 ;
      RECT   0.635000 143.675000   0.805000 143.845000 ;
      RECT   0.635000 144.895000   0.805000 145.065000 ;
      RECT   0.635000 146.115000   0.805000 146.285000 ;
      RECT   0.635000 147.335000   0.805000 147.505000 ;
      RECT   0.635000 148.555000   0.805000 148.725000 ;
      RECT   0.635000 149.775000   0.805000 149.945000 ;
      RECT   0.635000 150.995000   0.805000 151.165000 ;
      RECT   0.635000 152.215000   0.805000 152.385000 ;
      RECT   0.635000 153.435000   0.805000 153.605000 ;
      RECT   0.635000 154.655000   0.805000 154.825000 ;
      RECT   0.850000 156.415000   1.020000 156.585000 ;
      RECT   0.920000  -8.145000   1.090000  -7.975000 ;
      RECT   1.115000  -6.385000   1.285000  -6.215000 ;
      RECT   1.115000  -5.165000   1.285000  -4.995000 ;
      RECT   1.115000  -3.945000   1.285000  -3.775000 ;
      RECT   1.115000  -2.725000   1.285000  -2.555000 ;
      RECT   1.115000  -1.505000   1.285000  -1.335000 ;
      RECT   1.115000  -0.285000   1.285000  -0.115000 ;
      RECT   1.115000   0.935000   1.285000   1.105000 ;
      RECT   1.115000   2.155000   1.285000   2.325000 ;
      RECT   1.115000   3.375000   1.285000   3.545000 ;
      RECT   1.115000   4.595000   1.285000   4.765000 ;
      RECT   1.115000   5.815000   1.285000   5.985000 ;
      RECT   1.115000   7.035000   1.285000   7.205000 ;
      RECT   1.115000   8.255000   1.285000   8.425000 ;
      RECT   1.115000   9.475000   1.285000   9.645000 ;
      RECT   1.115000  10.695000   1.285000  10.865000 ;
      RECT   1.115000  11.915000   1.285000  12.085000 ;
      RECT   1.115000  13.135000   1.285000  13.305000 ;
      RECT   1.115000  14.355000   1.285000  14.525000 ;
      RECT   1.115000  15.575000   1.285000  15.745000 ;
      RECT   1.115000  16.795000   1.285000  16.965000 ;
      RECT   1.115000  18.015000   1.285000  18.185000 ;
      RECT   1.115000  19.235000   1.285000  19.405000 ;
      RECT   1.115000  20.455000   1.285000  20.625000 ;
      RECT   1.115000  21.675000   1.285000  21.845000 ;
      RECT   1.115000  22.895000   1.285000  23.065000 ;
      RECT   1.115000  24.115000   1.285000  24.285000 ;
      RECT   1.115000  25.335000   1.285000  25.505000 ;
      RECT   1.115000  26.555000   1.285000  26.725000 ;
      RECT   1.115000  27.775000   1.285000  27.945000 ;
      RECT   1.115000  28.995000   1.285000  29.165000 ;
      RECT   1.115000  30.215000   1.285000  30.385000 ;
      RECT   1.115000  31.435000   1.285000  31.605000 ;
      RECT   1.115000  32.655000   1.285000  32.825000 ;
      RECT   1.115000  33.875000   1.285000  34.045000 ;
      RECT   1.115000  35.095000   1.285000  35.265000 ;
      RECT   1.115000  36.315000   1.285000  36.485000 ;
      RECT   1.115000  37.535000   1.285000  37.705000 ;
      RECT   1.115000  38.755000   1.285000  38.925000 ;
      RECT   1.115000  39.975000   1.285000  40.145000 ;
      RECT   1.115000  41.195000   1.285000  41.365000 ;
      RECT   1.115000  42.415000   1.285000  42.585000 ;
      RECT   1.115000  43.635000   1.285000  43.805000 ;
      RECT   1.115000  44.855000   1.285000  45.025000 ;
      RECT   1.115000  46.075000   1.285000  46.245000 ;
      RECT   1.115000  47.295000   1.285000  47.465000 ;
      RECT   1.115000  48.515000   1.285000  48.685000 ;
      RECT   1.115000  49.735000   1.285000  49.905000 ;
      RECT   1.115000  50.955000   1.285000  51.125000 ;
      RECT   1.115000  52.175000   1.285000  52.345000 ;
      RECT   1.115000  53.395000   1.285000  53.565000 ;
      RECT   1.115000  54.615000   1.285000  54.785000 ;
      RECT   1.115000  55.835000   1.285000  56.005000 ;
      RECT   1.115000  57.055000   1.285000  57.225000 ;
      RECT   1.115000  58.275000   1.285000  58.445000 ;
      RECT   1.115000  59.495000   1.285000  59.665000 ;
      RECT   1.115000  60.715000   1.285000  60.885000 ;
      RECT   1.115000  61.935000   1.285000  62.105000 ;
      RECT   1.115000  63.155000   1.285000  63.325000 ;
      RECT   1.115000  64.375000   1.285000  64.545000 ;
      RECT   1.115000  65.595000   1.285000  65.765000 ;
      RECT   1.115000  66.815000   1.285000  66.985000 ;
      RECT   1.115000  68.035000   1.285000  68.205000 ;
      RECT   1.115000  69.255000   1.285000  69.425000 ;
      RECT   1.115000  70.475000   1.285000  70.645000 ;
      RECT   1.115000  71.695000   1.285000  71.865000 ;
      RECT   1.115000  72.915000   1.285000  73.085000 ;
      RECT   1.115000  74.135000   1.285000  74.305000 ;
      RECT   1.115000  75.355000   1.285000  75.525000 ;
      RECT   1.115000  76.575000   1.285000  76.745000 ;
      RECT   1.115000  77.795000   1.285000  77.965000 ;
      RECT   1.115000  79.015000   1.285000  79.185000 ;
      RECT   1.115000  80.235000   1.285000  80.405000 ;
      RECT   1.115000  81.455000   1.285000  81.625000 ;
      RECT   1.115000  82.675000   1.285000  82.845000 ;
      RECT   1.115000  83.895000   1.285000  84.065000 ;
      RECT   1.115000  85.115000   1.285000  85.285000 ;
      RECT   1.115000  86.335000   1.285000  86.505000 ;
      RECT   1.115000  87.555000   1.285000  87.725000 ;
      RECT   1.115000  88.775000   1.285000  88.945000 ;
      RECT   1.115000  89.995000   1.285000  90.165000 ;
      RECT   1.115000  91.215000   1.285000  91.385000 ;
      RECT   1.115000  92.435000   1.285000  92.605000 ;
      RECT   1.115000  93.655000   1.285000  93.825000 ;
      RECT   1.115000  94.875000   1.285000  95.045000 ;
      RECT   1.115000  96.095000   1.285000  96.265000 ;
      RECT   1.115000  97.315000   1.285000  97.485000 ;
      RECT   1.115000  98.535000   1.285000  98.705000 ;
      RECT   1.115000  99.755000   1.285000  99.925000 ;
      RECT   1.115000 100.975000   1.285000 101.145000 ;
      RECT   1.115000 102.195000   1.285000 102.365000 ;
      RECT   1.115000 103.415000   1.285000 103.585000 ;
      RECT   1.115000 104.635000   1.285000 104.805000 ;
      RECT   1.115000 105.855000   1.285000 106.025000 ;
      RECT   1.115000 107.075000   1.285000 107.245000 ;
      RECT   1.115000 108.295000   1.285000 108.465000 ;
      RECT   1.115000 109.515000   1.285000 109.685000 ;
      RECT   1.115000 110.735000   1.285000 110.905000 ;
      RECT   1.115000 111.955000   1.285000 112.125000 ;
      RECT   1.115000 113.175000   1.285000 113.345000 ;
      RECT   1.115000 114.395000   1.285000 114.565000 ;
      RECT   1.115000 115.615000   1.285000 115.785000 ;
      RECT   1.115000 116.835000   1.285000 117.005000 ;
      RECT   1.115000 118.055000   1.285000 118.225000 ;
      RECT   1.115000 119.275000   1.285000 119.445000 ;
      RECT   1.115000 120.495000   1.285000 120.665000 ;
      RECT   1.115000 121.715000   1.285000 121.885000 ;
      RECT   1.115000 122.935000   1.285000 123.105000 ;
      RECT   1.115000 124.155000   1.285000 124.325000 ;
      RECT   1.115000 125.375000   1.285000 125.545000 ;
      RECT   1.115000 126.595000   1.285000 126.765000 ;
      RECT   1.115000 127.815000   1.285000 127.985000 ;
      RECT   1.115000 129.035000   1.285000 129.205000 ;
      RECT   1.115000 130.255000   1.285000 130.425000 ;
      RECT   1.115000 131.475000   1.285000 131.645000 ;
      RECT   1.115000 132.695000   1.285000 132.865000 ;
      RECT   1.115000 133.915000   1.285000 134.085000 ;
      RECT   1.115000 135.135000   1.285000 135.305000 ;
      RECT   1.115000 136.355000   1.285000 136.525000 ;
      RECT   1.115000 137.575000   1.285000 137.745000 ;
      RECT   1.115000 138.795000   1.285000 138.965000 ;
      RECT   1.115000 140.015000   1.285000 140.185000 ;
      RECT   1.115000 141.235000   1.285000 141.405000 ;
      RECT   1.115000 142.455000   1.285000 142.625000 ;
      RECT   1.115000 143.675000   1.285000 143.845000 ;
      RECT   1.115000 144.895000   1.285000 145.065000 ;
      RECT   1.115000 146.115000   1.285000 146.285000 ;
      RECT   1.115000 147.335000   1.285000 147.505000 ;
      RECT   1.115000 148.555000   1.285000 148.725000 ;
      RECT   1.115000 149.775000   1.285000 149.945000 ;
      RECT   1.115000 150.995000   1.285000 151.165000 ;
      RECT   1.115000 152.215000   1.285000 152.385000 ;
      RECT   1.115000 153.435000   1.285000 153.605000 ;
      RECT   1.115000 154.655000   1.285000 154.825000 ;
      RECT   1.210000 156.415000   1.380000 156.585000 ;
      RECT   1.285000  -8.145000   1.455000  -7.975000 ;
      RECT   1.570000 156.415000   1.740000 156.585000 ;
      RECT   1.595000  -6.385000   1.765000  -6.215000 ;
      RECT   1.595000  -5.165000   1.765000  -4.995000 ;
      RECT   1.595000  -3.945000   1.765000  -3.775000 ;
      RECT   1.595000  -2.725000   1.765000  -2.555000 ;
      RECT   1.595000  -1.505000   1.765000  -1.335000 ;
      RECT   1.595000  -0.285000   1.765000  -0.115000 ;
      RECT   1.595000   0.935000   1.765000   1.105000 ;
      RECT   1.595000   2.155000   1.765000   2.325000 ;
      RECT   1.595000   3.375000   1.765000   3.545000 ;
      RECT   1.595000   4.595000   1.765000   4.765000 ;
      RECT   1.595000   5.815000   1.765000   5.985000 ;
      RECT   1.595000   7.035000   1.765000   7.205000 ;
      RECT   1.595000   8.255000   1.765000   8.425000 ;
      RECT   1.595000   9.475000   1.765000   9.645000 ;
      RECT   1.595000  10.695000   1.765000  10.865000 ;
      RECT   1.595000  11.915000   1.765000  12.085000 ;
      RECT   1.595000  13.135000   1.765000  13.305000 ;
      RECT   1.595000  14.355000   1.765000  14.525000 ;
      RECT   1.595000  15.575000   1.765000  15.745000 ;
      RECT   1.595000  16.795000   1.765000  16.965000 ;
      RECT   1.595000  18.015000   1.765000  18.185000 ;
      RECT   1.595000  19.235000   1.765000  19.405000 ;
      RECT   1.595000  20.455000   1.765000  20.625000 ;
      RECT   1.595000  21.675000   1.765000  21.845000 ;
      RECT   1.595000  22.895000   1.765000  23.065000 ;
      RECT   1.595000  24.115000   1.765000  24.285000 ;
      RECT   1.595000  25.335000   1.765000  25.505000 ;
      RECT   1.595000  26.555000   1.765000  26.725000 ;
      RECT   1.595000  27.775000   1.765000  27.945000 ;
      RECT   1.595000  28.995000   1.765000  29.165000 ;
      RECT   1.595000  30.215000   1.765000  30.385000 ;
      RECT   1.595000  31.435000   1.765000  31.605000 ;
      RECT   1.595000  32.655000   1.765000  32.825000 ;
      RECT   1.595000  33.875000   1.765000  34.045000 ;
      RECT   1.595000  35.095000   1.765000  35.265000 ;
      RECT   1.595000  36.315000   1.765000  36.485000 ;
      RECT   1.595000  37.535000   1.765000  37.705000 ;
      RECT   1.595000  38.755000   1.765000  38.925000 ;
      RECT   1.595000  39.975000   1.765000  40.145000 ;
      RECT   1.595000  41.195000   1.765000  41.365000 ;
      RECT   1.595000  42.415000   1.765000  42.585000 ;
      RECT   1.595000  43.635000   1.765000  43.805000 ;
      RECT   1.595000  44.855000   1.765000  45.025000 ;
      RECT   1.595000  46.075000   1.765000  46.245000 ;
      RECT   1.595000  47.295000   1.765000  47.465000 ;
      RECT   1.595000  48.515000   1.765000  48.685000 ;
      RECT   1.595000  49.735000   1.765000  49.905000 ;
      RECT   1.595000  50.955000   1.765000  51.125000 ;
      RECT   1.595000  52.175000   1.765000  52.345000 ;
      RECT   1.595000  53.395000   1.765000  53.565000 ;
      RECT   1.595000  54.615000   1.765000  54.785000 ;
      RECT   1.595000  55.835000   1.765000  56.005000 ;
      RECT   1.595000  57.055000   1.765000  57.225000 ;
      RECT   1.595000  58.275000   1.765000  58.445000 ;
      RECT   1.595000  59.495000   1.765000  59.665000 ;
      RECT   1.595000  60.715000   1.765000  60.885000 ;
      RECT   1.595000  61.935000   1.765000  62.105000 ;
      RECT   1.595000  63.155000   1.765000  63.325000 ;
      RECT   1.595000  64.375000   1.765000  64.545000 ;
      RECT   1.595000  65.595000   1.765000  65.765000 ;
      RECT   1.595000  66.815000   1.765000  66.985000 ;
      RECT   1.595000  68.035000   1.765000  68.205000 ;
      RECT   1.595000  69.255000   1.765000  69.425000 ;
      RECT   1.595000  70.475000   1.765000  70.645000 ;
      RECT   1.595000  71.695000   1.765000  71.865000 ;
      RECT   1.595000  72.915000   1.765000  73.085000 ;
      RECT   1.595000  74.135000   1.765000  74.305000 ;
      RECT   1.595000  75.355000   1.765000  75.525000 ;
      RECT   1.595000  76.575000   1.765000  76.745000 ;
      RECT   1.595000  77.795000   1.765000  77.965000 ;
      RECT   1.595000  79.015000   1.765000  79.185000 ;
      RECT   1.595000  80.235000   1.765000  80.405000 ;
      RECT   1.595000  81.455000   1.765000  81.625000 ;
      RECT   1.595000  82.675000   1.765000  82.845000 ;
      RECT   1.595000  83.895000   1.765000  84.065000 ;
      RECT   1.595000  85.115000   1.765000  85.285000 ;
      RECT   1.595000  86.335000   1.765000  86.505000 ;
      RECT   1.595000  87.555000   1.765000  87.725000 ;
      RECT   1.595000  88.775000   1.765000  88.945000 ;
      RECT   1.595000  89.995000   1.765000  90.165000 ;
      RECT   1.595000  91.215000   1.765000  91.385000 ;
      RECT   1.595000  92.435000   1.765000  92.605000 ;
      RECT   1.595000  93.655000   1.765000  93.825000 ;
      RECT   1.595000  94.875000   1.765000  95.045000 ;
      RECT   1.595000  96.095000   1.765000  96.265000 ;
      RECT   1.595000  97.315000   1.765000  97.485000 ;
      RECT   1.595000  98.535000   1.765000  98.705000 ;
      RECT   1.595000  99.755000   1.765000  99.925000 ;
      RECT   1.595000 100.975000   1.765000 101.145000 ;
      RECT   1.595000 102.195000   1.765000 102.365000 ;
      RECT   1.595000 103.415000   1.765000 103.585000 ;
      RECT   1.595000 104.635000   1.765000 104.805000 ;
      RECT   1.595000 105.855000   1.765000 106.025000 ;
      RECT   1.595000 107.075000   1.765000 107.245000 ;
      RECT   1.595000 108.295000   1.765000 108.465000 ;
      RECT   1.595000 109.515000   1.765000 109.685000 ;
      RECT   1.595000 110.735000   1.765000 110.905000 ;
      RECT   1.595000 111.955000   1.765000 112.125000 ;
      RECT   1.595000 113.175000   1.765000 113.345000 ;
      RECT   1.595000 114.395000   1.765000 114.565000 ;
      RECT   1.595000 115.615000   1.765000 115.785000 ;
      RECT   1.595000 116.835000   1.765000 117.005000 ;
      RECT   1.595000 118.055000   1.765000 118.225000 ;
      RECT   1.595000 119.275000   1.765000 119.445000 ;
      RECT   1.595000 120.495000   1.765000 120.665000 ;
      RECT   1.595000 121.715000   1.765000 121.885000 ;
      RECT   1.595000 122.935000   1.765000 123.105000 ;
      RECT   1.595000 124.155000   1.765000 124.325000 ;
      RECT   1.595000 125.375000   1.765000 125.545000 ;
      RECT   1.595000 126.595000   1.765000 126.765000 ;
      RECT   1.595000 127.815000   1.765000 127.985000 ;
      RECT   1.595000 129.035000   1.765000 129.205000 ;
      RECT   1.595000 130.255000   1.765000 130.425000 ;
      RECT   1.595000 131.475000   1.765000 131.645000 ;
      RECT   1.595000 132.695000   1.765000 132.865000 ;
      RECT   1.595000 133.915000   1.765000 134.085000 ;
      RECT   1.595000 135.135000   1.765000 135.305000 ;
      RECT   1.595000 136.355000   1.765000 136.525000 ;
      RECT   1.595000 137.575000   1.765000 137.745000 ;
      RECT   1.595000 138.795000   1.765000 138.965000 ;
      RECT   1.595000 140.015000   1.765000 140.185000 ;
      RECT   1.595000 141.235000   1.765000 141.405000 ;
      RECT   1.595000 142.455000   1.765000 142.625000 ;
      RECT   1.595000 143.675000   1.765000 143.845000 ;
      RECT   1.595000 144.895000   1.765000 145.065000 ;
      RECT   1.595000 146.115000   1.765000 146.285000 ;
      RECT   1.595000 147.335000   1.765000 147.505000 ;
      RECT   1.595000 148.555000   1.765000 148.725000 ;
      RECT   1.595000 149.775000   1.765000 149.945000 ;
      RECT   1.595000 150.995000   1.765000 151.165000 ;
      RECT   1.595000 152.215000   1.765000 152.385000 ;
      RECT   1.595000 153.435000   1.765000 153.605000 ;
      RECT   1.595000 154.655000   1.765000 154.825000 ;
      RECT   1.650000  -8.145000   1.820000  -7.975000 ;
      RECT   1.930000 156.415000   2.100000 156.585000 ;
      RECT   2.015000  -8.145000   2.185000  -7.975000 ;
      RECT   2.075000  -6.385000   2.245000  -6.215000 ;
      RECT   2.075000  -5.165000   2.245000  -4.995000 ;
      RECT   2.075000  -3.945000   2.245000  -3.775000 ;
      RECT   2.075000  -2.725000   2.245000  -2.555000 ;
      RECT   2.075000  -1.505000   2.245000  -1.335000 ;
      RECT   2.075000  -0.285000   2.245000  -0.115000 ;
      RECT   2.075000   0.935000   2.245000   1.105000 ;
      RECT   2.075000   2.155000   2.245000   2.325000 ;
      RECT   2.075000   3.375000   2.245000   3.545000 ;
      RECT   2.075000   4.595000   2.245000   4.765000 ;
      RECT   2.075000   5.815000   2.245000   5.985000 ;
      RECT   2.075000   7.035000   2.245000   7.205000 ;
      RECT   2.075000   8.255000   2.245000   8.425000 ;
      RECT   2.075000   9.475000   2.245000   9.645000 ;
      RECT   2.075000  10.695000   2.245000  10.865000 ;
      RECT   2.075000  11.915000   2.245000  12.085000 ;
      RECT   2.075000  13.135000   2.245000  13.305000 ;
      RECT   2.075000  14.355000   2.245000  14.525000 ;
      RECT   2.075000  15.575000   2.245000  15.745000 ;
      RECT   2.075000  16.795000   2.245000  16.965000 ;
      RECT   2.075000  18.015000   2.245000  18.185000 ;
      RECT   2.075000  19.235000   2.245000  19.405000 ;
      RECT   2.075000  20.455000   2.245000  20.625000 ;
      RECT   2.075000  21.675000   2.245000  21.845000 ;
      RECT   2.075000  22.895000   2.245000  23.065000 ;
      RECT   2.075000  24.115000   2.245000  24.285000 ;
      RECT   2.075000  25.335000   2.245000  25.505000 ;
      RECT   2.075000  26.555000   2.245000  26.725000 ;
      RECT   2.075000  27.775000   2.245000  27.945000 ;
      RECT   2.075000  28.995000   2.245000  29.165000 ;
      RECT   2.075000  30.215000   2.245000  30.385000 ;
      RECT   2.075000  31.435000   2.245000  31.605000 ;
      RECT   2.075000  32.655000   2.245000  32.825000 ;
      RECT   2.075000  33.875000   2.245000  34.045000 ;
      RECT   2.075000  35.095000   2.245000  35.265000 ;
      RECT   2.075000  36.315000   2.245000  36.485000 ;
      RECT   2.075000  37.535000   2.245000  37.705000 ;
      RECT   2.075000  38.755000   2.245000  38.925000 ;
      RECT   2.075000  39.975000   2.245000  40.145000 ;
      RECT   2.075000  41.195000   2.245000  41.365000 ;
      RECT   2.075000  42.415000   2.245000  42.585000 ;
      RECT   2.075000  43.635000   2.245000  43.805000 ;
      RECT   2.075000  44.855000   2.245000  45.025000 ;
      RECT   2.075000  46.075000   2.245000  46.245000 ;
      RECT   2.075000  47.295000   2.245000  47.465000 ;
      RECT   2.075000  48.515000   2.245000  48.685000 ;
      RECT   2.075000  49.735000   2.245000  49.905000 ;
      RECT   2.075000  50.955000   2.245000  51.125000 ;
      RECT   2.075000  52.175000   2.245000  52.345000 ;
      RECT   2.075000  53.395000   2.245000  53.565000 ;
      RECT   2.075000  54.615000   2.245000  54.785000 ;
      RECT   2.075000  55.835000   2.245000  56.005000 ;
      RECT   2.075000  57.055000   2.245000  57.225000 ;
      RECT   2.075000  58.275000   2.245000  58.445000 ;
      RECT   2.075000  59.495000   2.245000  59.665000 ;
      RECT   2.075000  60.715000   2.245000  60.885000 ;
      RECT   2.075000  61.935000   2.245000  62.105000 ;
      RECT   2.075000  63.155000   2.245000  63.325000 ;
      RECT   2.075000  64.375000   2.245000  64.545000 ;
      RECT   2.075000  65.595000   2.245000  65.765000 ;
      RECT   2.075000  66.815000   2.245000  66.985000 ;
      RECT   2.075000  68.035000   2.245000  68.205000 ;
      RECT   2.075000  69.255000   2.245000  69.425000 ;
      RECT   2.075000  70.475000   2.245000  70.645000 ;
      RECT   2.075000  71.695000   2.245000  71.865000 ;
      RECT   2.075000  72.915000   2.245000  73.085000 ;
      RECT   2.075000  74.135000   2.245000  74.305000 ;
      RECT   2.075000  75.355000   2.245000  75.525000 ;
      RECT   2.075000  76.575000   2.245000  76.745000 ;
      RECT   2.075000  77.795000   2.245000  77.965000 ;
      RECT   2.075000  79.015000   2.245000  79.185000 ;
      RECT   2.075000  80.235000   2.245000  80.405000 ;
      RECT   2.075000  81.455000   2.245000  81.625000 ;
      RECT   2.075000  82.675000   2.245000  82.845000 ;
      RECT   2.075000  83.895000   2.245000  84.065000 ;
      RECT   2.075000  85.115000   2.245000  85.285000 ;
      RECT   2.075000  86.335000   2.245000  86.505000 ;
      RECT   2.075000  87.555000   2.245000  87.725000 ;
      RECT   2.075000  88.775000   2.245000  88.945000 ;
      RECT   2.075000  89.995000   2.245000  90.165000 ;
      RECT   2.075000  91.215000   2.245000  91.385000 ;
      RECT   2.075000  92.435000   2.245000  92.605000 ;
      RECT   2.075000  93.655000   2.245000  93.825000 ;
      RECT   2.075000  94.875000   2.245000  95.045000 ;
      RECT   2.075000  96.095000   2.245000  96.265000 ;
      RECT   2.075000  97.315000   2.245000  97.485000 ;
      RECT   2.075000  98.535000   2.245000  98.705000 ;
      RECT   2.075000  99.755000   2.245000  99.925000 ;
      RECT   2.075000 100.975000   2.245000 101.145000 ;
      RECT   2.075000 102.195000   2.245000 102.365000 ;
      RECT   2.075000 103.415000   2.245000 103.585000 ;
      RECT   2.075000 104.635000   2.245000 104.805000 ;
      RECT   2.075000 105.855000   2.245000 106.025000 ;
      RECT   2.075000 107.075000   2.245000 107.245000 ;
      RECT   2.075000 108.295000   2.245000 108.465000 ;
      RECT   2.075000 109.515000   2.245000 109.685000 ;
      RECT   2.075000 110.735000   2.245000 110.905000 ;
      RECT   2.075000 111.955000   2.245000 112.125000 ;
      RECT   2.075000 113.175000   2.245000 113.345000 ;
      RECT   2.075000 114.395000   2.245000 114.565000 ;
      RECT   2.075000 115.615000   2.245000 115.785000 ;
      RECT   2.075000 116.835000   2.245000 117.005000 ;
      RECT   2.075000 118.055000   2.245000 118.225000 ;
      RECT   2.075000 119.275000   2.245000 119.445000 ;
      RECT   2.075000 120.495000   2.245000 120.665000 ;
      RECT   2.075000 121.715000   2.245000 121.885000 ;
      RECT   2.075000 122.935000   2.245000 123.105000 ;
      RECT   2.075000 124.155000   2.245000 124.325000 ;
      RECT   2.075000 125.375000   2.245000 125.545000 ;
      RECT   2.075000 126.595000   2.245000 126.765000 ;
      RECT   2.075000 127.815000   2.245000 127.985000 ;
      RECT   2.075000 129.035000   2.245000 129.205000 ;
      RECT   2.075000 130.255000   2.245000 130.425000 ;
      RECT   2.075000 131.475000   2.245000 131.645000 ;
      RECT   2.075000 132.695000   2.245000 132.865000 ;
      RECT   2.075000 133.915000   2.245000 134.085000 ;
      RECT   2.075000 135.135000   2.245000 135.305000 ;
      RECT   2.075000 136.355000   2.245000 136.525000 ;
      RECT   2.075000 137.575000   2.245000 137.745000 ;
      RECT   2.075000 138.795000   2.245000 138.965000 ;
      RECT   2.075000 140.015000   2.245000 140.185000 ;
      RECT   2.075000 141.235000   2.245000 141.405000 ;
      RECT   2.075000 142.455000   2.245000 142.625000 ;
      RECT   2.075000 143.675000   2.245000 143.845000 ;
      RECT   2.075000 144.895000   2.245000 145.065000 ;
      RECT   2.075000 146.115000   2.245000 146.285000 ;
      RECT   2.075000 147.335000   2.245000 147.505000 ;
      RECT   2.075000 148.555000   2.245000 148.725000 ;
      RECT   2.075000 149.775000   2.245000 149.945000 ;
      RECT   2.075000 150.995000   2.245000 151.165000 ;
      RECT   2.075000 152.215000   2.245000 152.385000 ;
      RECT   2.075000 153.435000   2.245000 153.605000 ;
      RECT   2.075000 154.655000   2.245000 154.825000 ;
      RECT   2.290000 156.415000   2.460000 156.585000 ;
      RECT   2.380000  -8.145000   2.550000  -7.975000 ;
      RECT   2.650000 156.415000   2.820000 156.585000 ;
      RECT   2.745000  -8.145000   2.915000  -7.975000 ;
      RECT   3.010000 156.415000   3.180000 156.585000 ;
      RECT   3.110000  -8.145000   3.280000  -7.975000 ;
      RECT   3.370000 156.415000   3.540000 156.585000 ;
      RECT   3.475000  -8.145000   3.645000  -7.975000 ;
      RECT   3.730000 156.415000   3.900000 156.585000 ;
      RECT   3.840000  -8.145000   4.010000  -7.975000 ;
      RECT   4.090000 156.415000   4.260000 156.585000 ;
      RECT   4.205000  -8.145000   4.375000  -7.975000 ;
      RECT   4.450000 156.415000   4.620000 156.585000 ;
      RECT   4.570000  -8.145000   4.740000  -7.975000 ;
      RECT   4.810000 156.415000   4.980000 156.585000 ;
      RECT   4.935000  -8.145000   5.105000  -7.975000 ;
      RECT   5.170000 156.415000   5.340000 156.585000 ;
      RECT   5.300000  -8.145000   5.470000  -7.975000 ;
      RECT   5.530000 156.415000   5.700000 156.585000 ;
      RECT   5.665000  -8.145000   5.835000  -7.975000 ;
      RECT   5.890000 156.415000   6.060000 156.585000 ;
      RECT   6.030000  -8.145000   6.200000  -7.975000 ;
      RECT   6.250000 156.415000   6.420000 156.585000 ;
      RECT   6.395000  -8.145000   6.565000  -7.975000 ;
      RECT   6.610000 156.415000   6.780000 156.585000 ;
      RECT   6.760000  -8.145000   6.930000  -7.975000 ;
      RECT   6.970000 156.415000   7.140000 156.585000 ;
      RECT   7.125000  -8.145000   7.295000  -7.975000 ;
      RECT   7.330000 156.415000   7.500000 156.585000 ;
      RECT   7.490000  -8.145000   7.660000  -7.975000 ;
      RECT   7.690000 156.415000   7.860000 156.585000 ;
      RECT   7.855000  -8.145000   8.025000  -7.975000 ;
      RECT   8.050000 156.415000   8.220000 156.585000 ;
      RECT   8.220000  -8.145000   8.390000  -7.975000 ;
      RECT   8.410000 156.415000   8.580000 156.585000 ;
      RECT   8.585000  -8.145000   8.755000  -7.975000 ;
      RECT   8.770000 156.415000   8.940000 156.585000 ;
      RECT   8.950000  -8.145000   9.120000  -7.975000 ;
      RECT   9.130000 156.415000   9.300000 156.585000 ;
      RECT   9.315000  -8.145000   9.485000  -7.975000 ;
      RECT   9.490000 156.415000   9.660000 156.585000 ;
      RECT   9.680000  -8.145000   9.850000  -7.975000 ;
      RECT   9.850000 156.415000  10.020000 156.585000 ;
      RECT  10.045000  -8.145000  10.215000  -7.975000 ;
      RECT  10.210000 156.415000  10.380000 156.585000 ;
      RECT  10.410000  -8.145000  10.580000  -7.975000 ;
      RECT  10.570000 156.415000  10.740000 156.585000 ;
      RECT  10.775000  -8.145000  10.945000  -7.975000 ;
      RECT  10.930000 156.415000  11.100000 156.585000 ;
      RECT  11.140000  -8.145000  11.310000  -7.975000 ;
      RECT  11.290000 156.415000  11.460000 156.585000 ;
      RECT  11.505000  -8.145000  11.675000  -7.975000 ;
      RECT  11.650000 156.415000  11.820000 156.585000 ;
      RECT  11.870000  -8.145000  12.040000  -7.975000 ;
      RECT  12.010000 156.415000  12.180000 156.585000 ;
      RECT  12.235000  -8.145000  12.405000  -7.975000 ;
      RECT  12.370000 156.415000  12.540000 156.585000 ;
      RECT  12.600000  -8.145000  12.770000  -7.975000 ;
      RECT  12.730000 156.415000  12.900000 156.585000 ;
      RECT  12.965000  -8.145000  13.135000  -7.975000 ;
      RECT  13.090000 156.415000  13.260000 156.585000 ;
      RECT  13.330000  -8.145000  13.500000  -7.975000 ;
      RECT  13.450000 156.415000  13.620000 156.585000 ;
      RECT  13.695000  -8.145000  13.865000  -7.975000 ;
      RECT  13.810000 156.415000  13.980000 156.585000 ;
      RECT  14.060000  -8.145000  14.230000  -7.975000 ;
      RECT  14.170000 156.415000  14.340000 156.585000 ;
      RECT  14.425000  -8.145000  14.595000  -7.975000 ;
      RECT  14.530000 156.415000  14.700000 156.585000 ;
      RECT  14.790000  -8.145000  14.960000  -7.975000 ;
      RECT  14.890000 156.415000  15.060000 156.585000 ;
      RECT  15.155000  -8.145000  15.325000  -7.975000 ;
      RECT  15.250000 156.415000  15.420000 156.585000 ;
      RECT  15.520000  -8.145000  15.690000  -7.975000 ;
      RECT  15.610000 156.415000  15.780000 156.585000 ;
      RECT  15.885000  -8.145000  16.055000  -7.975000 ;
      RECT  15.970000 156.415000  16.140000 156.585000 ;
      RECT  16.250000  -8.145000  16.420000  -7.975000 ;
      RECT  16.330000 156.415000  16.500000 156.585000 ;
      RECT  16.615000  -8.145000  16.785000  -7.975000 ;
      RECT  16.690000 156.415000  16.860000 156.585000 ;
      RECT  16.980000  -8.145000  17.150000  -7.975000 ;
      RECT  17.050000 156.415000  17.220000 156.585000 ;
      RECT  17.340000  -8.145000  17.510000  -7.975000 ;
      RECT  17.410000 156.415000  17.580000 156.585000 ;
      RECT  17.700000  -8.145000  17.870000  -7.975000 ;
      RECT  17.770000 156.415000  17.940000 156.585000 ;
      RECT  18.060000  -8.145000  18.230000  -7.975000 ;
      RECT  18.130000 156.415000  18.300000 156.585000 ;
      RECT  18.420000  -8.145000  18.590000  -7.975000 ;
      RECT  18.490000 156.415000  18.660000 156.585000 ;
      RECT  18.780000  -8.145000  18.950000  -7.975000 ;
      RECT  18.850000 156.415000  19.020000 156.585000 ;
      RECT  19.140000  -8.145000  19.310000  -7.975000 ;
      RECT  19.210000 156.415000  19.380000 156.585000 ;
      RECT  19.500000  -8.145000  19.670000  -7.975000 ;
      RECT  19.570000 156.415000  19.740000 156.585000 ;
      RECT  19.860000  -8.145000  20.030000  -7.975000 ;
      RECT  19.930000 156.415000  20.100000 156.585000 ;
      RECT  20.220000  -8.145000  20.390000  -7.975000 ;
      RECT  20.290000 156.415000  20.460000 156.585000 ;
      RECT  20.580000  -8.145000  20.750000  -7.975000 ;
      RECT  20.650000 156.415000  20.820000 156.585000 ;
      RECT  20.940000  -8.145000  21.110000  -7.975000 ;
      RECT  21.010000 156.415000  21.180000 156.585000 ;
      RECT  21.300000  -8.145000  21.470000  -7.975000 ;
      RECT  21.370000 156.415000  21.540000 156.585000 ;
      RECT  21.660000  -8.145000  21.830000  -7.975000 ;
      RECT  21.730000 156.415000  21.900000 156.585000 ;
      RECT  22.020000  -8.145000  22.190000  -7.975000 ;
      RECT  22.090000 156.415000  22.260000 156.585000 ;
      RECT  22.380000  -8.145000  22.550000  -7.975000 ;
      RECT  22.450000 156.415000  22.620000 156.585000 ;
      RECT  22.740000  -8.145000  22.910000  -7.975000 ;
      RECT  22.810000 156.415000  22.980000 156.585000 ;
      RECT  23.100000  -8.145000  23.270000  -7.975000 ;
      RECT  23.170000 156.415000  23.340000 156.585000 ;
      RECT  23.460000  -8.145000  23.630000  -7.975000 ;
      RECT  23.530000 156.415000  23.700000 156.585000 ;
      RECT  23.820000  -8.145000  23.990000  -7.975000 ;
      RECT  23.890000 156.415000  24.060000 156.585000 ;
      RECT  24.180000  -8.145000  24.350000  -7.975000 ;
      RECT  24.250000 156.415000  24.420000 156.585000 ;
      RECT  24.540000  -8.145000  24.710000  -7.975000 ;
      RECT  24.610000 156.415000  24.780000 156.585000 ;
      RECT  24.900000  -8.145000  25.070000  -7.975000 ;
      RECT  24.970000 156.415000  25.140000 156.585000 ;
      RECT  25.260000  -8.145000  25.430000  -7.975000 ;
      RECT  25.330000 156.415000  25.500000 156.585000 ;
      RECT  25.620000  -8.145000  25.790000  -7.975000 ;
      RECT  25.690000 156.415000  25.860000 156.585000 ;
      RECT  25.980000  -8.145000  26.150000  -7.975000 ;
      RECT  26.050000 156.415000  26.220000 156.585000 ;
      RECT  26.340000  -8.145000  26.510000  -7.975000 ;
      RECT  26.410000 156.415000  26.580000 156.585000 ;
      RECT  26.700000  -8.145000  26.870000  -7.975000 ;
      RECT  26.770000 156.415000  26.940000 156.585000 ;
      RECT  27.060000  -8.145000  27.230000  -7.975000 ;
      RECT  27.130000 156.415000  27.300000 156.585000 ;
      RECT  27.420000  -8.145000  27.590000  -7.975000 ;
      RECT  27.490000 156.415000  27.660000 156.585000 ;
      RECT  27.780000  -8.145000  27.950000  -7.975000 ;
      RECT  27.850000 156.415000  28.020000 156.585000 ;
      RECT  28.140000  -8.145000  28.310000  -7.975000 ;
      RECT  28.210000 156.415000  28.380000 156.585000 ;
      RECT  28.500000  -8.145000  28.670000  -7.975000 ;
      RECT  28.570000 156.415000  28.740000 156.585000 ;
      RECT  28.860000  -8.145000  29.030000  -7.975000 ;
      RECT  28.930000 156.415000  29.100000 156.585000 ;
      RECT  29.220000  -8.145000  29.390000  -7.975000 ;
      RECT  29.290000 156.415000  29.460000 156.585000 ;
      RECT  29.580000  -8.145000  29.750000  -7.975000 ;
      RECT  29.650000 156.415000  29.820000 156.585000 ;
      RECT  29.940000  -8.145000  30.110000  -7.975000 ;
      RECT  30.010000 156.415000  30.180000 156.585000 ;
      RECT  30.300000  -8.145000  30.470000  -7.975000 ;
      RECT  30.370000 156.415000  30.540000 156.585000 ;
      RECT  30.660000  -8.145000  30.830000  -7.975000 ;
      RECT  30.730000 156.415000  30.900000 156.585000 ;
      RECT  31.020000  -8.145000  31.190000  -7.975000 ;
      RECT  31.090000 156.415000  31.260000 156.585000 ;
      RECT  31.380000  -8.145000  31.550000  -7.975000 ;
      RECT  31.450000 156.415000  31.620000 156.585000 ;
      RECT  31.740000  -8.145000  31.910000  -7.975000 ;
      RECT  31.810000 156.415000  31.980000 156.585000 ;
      RECT  32.100000  -8.145000  32.270000  -7.975000 ;
      RECT  32.170000 156.415000  32.340000 156.585000 ;
      RECT  32.460000  -8.145000  32.630000  -7.975000 ;
      RECT  32.530000 156.415000  32.700000 156.585000 ;
      RECT  32.820000  -8.145000  32.990000  -7.975000 ;
      RECT  32.890000 156.415000  33.060000 156.585000 ;
      RECT  33.180000  -8.145000  33.350000  -7.975000 ;
      RECT  33.250000 156.415000  33.420000 156.585000 ;
      RECT  33.540000  -8.145000  33.710000  -7.975000 ;
      RECT  33.610000 156.415000  33.780000 156.585000 ;
      RECT  33.900000  -8.145000  34.070000  -7.975000 ;
      RECT  33.970000 156.415000  34.140000 156.585000 ;
      RECT  34.260000  -8.145000  34.430000  -7.975000 ;
      RECT  34.330000 156.415000  34.500000 156.585000 ;
      RECT  34.620000  -8.145000  34.790000  -7.975000 ;
      RECT  34.690000 156.415000  34.860000 156.585000 ;
      RECT  34.980000  -8.145000  35.150000  -7.975000 ;
      RECT  35.050000 156.415000  35.220000 156.585000 ;
      RECT  35.340000  -8.145000  35.510000  -7.975000 ;
      RECT  35.410000 156.415000  35.580000 156.585000 ;
      RECT  35.700000  -8.145000  35.870000  -7.975000 ;
      RECT  35.770000 156.415000  35.940000 156.585000 ;
      RECT  36.060000  -8.145000  36.230000  -7.975000 ;
      RECT  36.130000 156.415000  36.300000 156.585000 ;
      RECT  36.420000  -8.145000  36.590000  -7.975000 ;
      RECT  36.490000 156.415000  36.660000 156.585000 ;
      RECT  36.780000  -8.145000  36.950000  -7.975000 ;
      RECT  36.850000 156.415000  37.020000 156.585000 ;
      RECT  37.140000  -8.145000  37.310000  -7.975000 ;
      RECT  37.210000 156.415000  37.380000 156.585000 ;
      RECT  37.500000  -8.145000  37.670000  -7.975000 ;
      RECT  37.570000 156.415000  37.740000 156.585000 ;
      RECT  37.860000  -8.145000  38.030000  -7.975000 ;
      RECT  37.930000 156.415000  38.100000 156.585000 ;
      RECT  38.220000  -8.145000  38.390000  -7.975000 ;
      RECT  38.290000 156.415000  38.460000 156.585000 ;
      RECT  38.580000  -8.145000  38.750000  -7.975000 ;
      RECT  38.650000 156.415000  38.820000 156.585000 ;
      RECT  38.940000  -8.145000  39.110000  -7.975000 ;
      RECT  39.010000 156.415000  39.180000 156.585000 ;
      RECT  39.300000  -8.145000  39.470000  -7.975000 ;
      RECT  39.370000 156.415000  39.540000 156.585000 ;
      RECT  39.660000  -8.145000  39.830000  -7.975000 ;
      RECT  39.730000 156.415000  39.900000 156.585000 ;
      RECT  40.020000  -8.145000  40.190000  -7.975000 ;
      RECT  40.090000 156.415000  40.260000 156.585000 ;
      RECT  40.380000  -8.145000  40.550000  -7.975000 ;
      RECT  40.450000 156.415000  40.620000 156.585000 ;
      RECT  40.740000  -8.145000  40.910000  -7.975000 ;
      RECT  40.810000 156.415000  40.980000 156.585000 ;
      RECT  41.100000  -8.145000  41.270000  -7.975000 ;
      RECT  41.170000 156.415000  41.340000 156.585000 ;
      RECT  41.460000  -8.145000  41.630000  -7.975000 ;
      RECT  41.530000 156.415000  41.700000 156.585000 ;
      RECT  41.820000  -8.145000  41.990000  -7.975000 ;
      RECT  41.890000 156.415000  42.060000 156.585000 ;
      RECT  42.180000  -8.145000  42.350000  -7.975000 ;
      RECT  42.250000 156.415000  42.420000 156.585000 ;
      RECT  42.540000  -8.145000  42.710000  -7.975000 ;
      RECT  42.610000 156.415000  42.780000 156.585000 ;
      RECT  42.900000  -8.145000  43.070000  -7.975000 ;
      RECT  42.970000 156.415000  43.140000 156.585000 ;
      RECT  43.260000  -8.145000  43.430000  -7.975000 ;
      RECT  43.330000 156.415000  43.500000 156.585000 ;
      RECT  43.620000  -8.145000  43.790000  -7.975000 ;
      RECT  43.690000 156.415000  43.860000 156.585000 ;
      RECT  43.980000  -8.145000  44.150000  -7.975000 ;
      RECT  44.050000 156.415000  44.220000 156.585000 ;
      RECT  44.340000  -8.145000  44.510000  -7.975000 ;
      RECT  44.410000 156.415000  44.580000 156.585000 ;
      RECT  44.700000  -8.145000  44.870000  -7.975000 ;
      RECT  44.770000 156.415000  44.940000 156.585000 ;
      RECT  45.060000  -8.145000  45.230000  -7.975000 ;
      RECT  45.130000 156.415000  45.300000 156.585000 ;
      RECT  45.420000  -8.145000  45.590000  -7.975000 ;
      RECT  45.490000 156.415000  45.660000 156.585000 ;
      RECT  45.780000  -8.145000  45.950000  -7.975000 ;
      RECT  45.850000 156.415000  46.020000 156.585000 ;
      RECT  46.140000  -8.145000  46.310000  -7.975000 ;
      RECT  46.210000 156.415000  46.380000 156.585000 ;
      RECT  46.500000  -8.145000  46.670000  -7.975000 ;
      RECT  46.570000 156.415000  46.740000 156.585000 ;
      RECT  46.860000  -8.145000  47.030000  -7.975000 ;
      RECT  46.930000 156.415000  47.100000 156.585000 ;
      RECT  47.220000  -8.145000  47.390000  -7.975000 ;
      RECT  47.290000 156.415000  47.460000 156.585000 ;
      RECT  47.580000  -8.145000  47.750000  -7.975000 ;
      RECT  47.650000 156.415000  47.820000 156.585000 ;
      RECT  47.940000  -8.145000  48.110000  -7.975000 ;
      RECT  48.010000 156.415000  48.180000 156.585000 ;
      RECT  48.300000  -8.145000  48.470000  -7.975000 ;
      RECT  48.370000 156.415000  48.540000 156.585000 ;
      RECT  48.660000  -8.145000  48.830000  -7.975000 ;
      RECT  48.730000 156.415000  48.900000 156.585000 ;
      RECT  49.020000  -8.145000  49.190000  -7.975000 ;
      RECT  49.090000 156.415000  49.260000 156.585000 ;
      RECT  49.380000  -8.145000  49.550000  -7.975000 ;
      RECT  49.450000 156.415000  49.620000 156.585000 ;
      RECT  49.740000  -8.145000  49.910000  -7.975000 ;
      RECT  49.810000 156.415000  49.980000 156.585000 ;
      RECT  50.100000  -8.145000  50.270000  -7.975000 ;
      RECT  50.170000 156.415000  50.340000 156.585000 ;
      RECT  50.460000  -8.145000  50.630000  -7.975000 ;
      RECT  50.530000 156.415000  50.700000 156.585000 ;
      RECT  50.820000  -8.145000  50.990000  -7.975000 ;
      RECT  50.890000 156.415000  51.060000 156.585000 ;
      RECT  51.180000  -8.145000  51.350000  -7.975000 ;
      RECT  51.250000 156.415000  51.420000 156.585000 ;
      RECT  51.540000  -8.145000  51.710000  -7.975000 ;
      RECT  51.610000 156.415000  51.780000 156.585000 ;
      RECT  51.900000  -8.145000  52.070000  -7.975000 ;
      RECT  51.970000 156.415000  52.140000 156.585000 ;
      RECT  52.260000  -8.145000  52.430000  -7.975000 ;
      RECT  52.330000 156.415000  52.500000 156.585000 ;
      RECT  52.620000  -8.145000  52.790000  -7.975000 ;
      RECT  52.690000 156.415000  52.860000 156.585000 ;
      RECT  52.980000  -8.145000  53.150000  -7.975000 ;
      RECT  53.050000 156.415000  53.220000 156.585000 ;
      RECT  53.340000  -8.145000  53.510000  -7.975000 ;
      RECT  53.410000 156.415000  53.580000 156.585000 ;
      RECT  53.700000  -8.145000  53.870000  -7.975000 ;
      RECT  53.770000 156.415000  53.940000 156.585000 ;
      RECT  54.060000  -8.145000  54.230000  -7.975000 ;
      RECT  54.130000 156.415000  54.300000 156.585000 ;
      RECT  54.420000  -8.145000  54.590000  -7.975000 ;
      RECT  54.490000 156.415000  54.660000 156.585000 ;
      RECT  54.780000  -8.145000  54.950000  -7.975000 ;
      RECT  54.850000 156.415000  55.020000 156.585000 ;
      RECT  55.140000  -8.145000  55.310000  -7.975000 ;
      RECT  55.210000 156.415000  55.380000 156.585000 ;
      RECT  55.500000  -8.145000  55.670000  -7.975000 ;
      RECT  55.570000 156.415000  55.740000 156.585000 ;
      RECT  55.860000  -8.145000  56.030000  -7.975000 ;
      RECT  55.930000 156.415000  56.100000 156.585000 ;
      RECT  56.220000  -8.145000  56.390000  -7.975000 ;
      RECT  56.290000 156.415000  56.460000 156.585000 ;
      RECT  56.580000  -8.145000  56.750000  -7.975000 ;
      RECT  56.650000 156.415000  56.820000 156.585000 ;
      RECT  56.940000  -8.145000  57.110000  -7.975000 ;
      RECT  57.010000 156.415000  57.180000 156.585000 ;
      RECT  57.300000  -8.145000  57.470000  -7.975000 ;
      RECT  57.370000 156.415000  57.540000 156.585000 ;
      RECT  57.660000  -8.145000  57.830000  -7.975000 ;
      RECT  57.730000 156.415000  57.900000 156.585000 ;
      RECT  58.020000  -8.145000  58.190000  -7.975000 ;
      RECT  58.090000 156.415000  58.260000 156.585000 ;
      RECT  58.380000  -8.145000  58.550000  -7.975000 ;
      RECT  58.450000 156.415000  58.620000 156.585000 ;
      RECT  58.740000  -8.145000  58.910000  -7.975000 ;
      RECT  58.810000 156.415000  58.980000 156.585000 ;
      RECT  59.100000  -8.145000  59.270000  -7.975000 ;
      RECT  59.170000 156.415000  59.340000 156.585000 ;
      RECT  59.460000  -8.145000  59.630000  -7.975000 ;
      RECT  59.530000 156.415000  59.700000 156.585000 ;
      RECT  59.820000  -8.145000  59.990000  -7.975000 ;
      RECT  59.890000 156.415000  60.060000 156.585000 ;
      RECT  60.180000  -8.145000  60.350000  -7.975000 ;
      RECT  60.250000 156.415000  60.420000 156.585000 ;
      RECT  60.540000  -8.145000  60.710000  -7.975000 ;
      RECT  60.610000 156.415000  60.780000 156.585000 ;
      RECT  60.900000  -8.145000  61.070000  -7.975000 ;
      RECT  60.970000 156.415000  61.140000 156.585000 ;
      RECT  61.260000  -8.145000  61.430000  -7.975000 ;
      RECT  61.330000 156.415000  61.500000 156.585000 ;
      RECT  61.620000  -8.145000  61.790000  -7.975000 ;
      RECT  61.690000 156.415000  61.860000 156.585000 ;
      RECT  61.980000  -8.145000  62.150000  -7.975000 ;
      RECT  62.050000 156.415000  62.220000 156.585000 ;
      RECT  62.340000  -8.145000  62.510000  -7.975000 ;
      RECT  62.410000 156.415000  62.580000 156.585000 ;
      RECT  62.700000  -8.145000  62.870000  -7.975000 ;
      RECT  62.770000 156.415000  62.940000 156.585000 ;
      RECT  63.060000  -8.145000  63.230000  -7.975000 ;
      RECT  63.130000 156.415000  63.300000 156.585000 ;
      RECT  63.420000  -8.145000  63.590000  -7.975000 ;
      RECT  63.490000 156.415000  63.660000 156.585000 ;
      RECT  63.780000  -8.145000  63.950000  -7.975000 ;
      RECT  63.850000 156.415000  64.020000 156.585000 ;
      RECT  64.140000  -8.145000  64.310000  -7.975000 ;
      RECT  64.210000 156.415000  64.380000 156.585000 ;
      RECT  64.500000  -8.145000  64.670000  -7.975000 ;
      RECT  64.570000 156.415000  64.740000 156.585000 ;
      RECT  64.860000  -8.145000  65.030000  -7.975000 ;
      RECT  64.930000 156.415000  65.100000 156.585000 ;
      RECT  65.220000  -8.145000  65.390000  -7.975000 ;
      RECT  65.290000 156.415000  65.460000 156.585000 ;
      RECT  65.580000  -8.145000  65.750000  -7.975000 ;
      RECT  65.650000 156.415000  65.820000 156.585000 ;
      RECT  65.940000  -8.145000  66.110000  -7.975000 ;
      RECT  66.010000 156.415000  66.180000 156.585000 ;
      RECT  66.300000  -8.145000  66.470000  -7.975000 ;
      RECT  66.370000 156.415000  66.540000 156.585000 ;
      RECT  66.660000  -8.145000  66.830000  -7.975000 ;
      RECT  66.730000 156.415000  66.900000 156.585000 ;
      RECT  67.020000  -8.145000  67.190000  -7.975000 ;
      RECT  67.090000 156.415000  67.260000 156.585000 ;
      RECT  67.380000  -8.145000  67.550000  -7.975000 ;
      RECT  67.450000 156.415000  67.620000 156.585000 ;
      RECT  67.740000  -8.145000  67.910000  -7.975000 ;
      RECT  67.810000 156.415000  67.980000 156.585000 ;
      RECT  68.100000  -8.145000  68.270000  -7.975000 ;
      RECT  68.170000 156.415000  68.340000 156.585000 ;
      RECT  68.460000  -8.145000  68.630000  -7.975000 ;
      RECT  68.530000 156.415000  68.700000 156.585000 ;
      RECT  68.820000  -8.145000  68.990000  -7.975000 ;
      RECT  68.890000 156.415000  69.060000 156.585000 ;
      RECT  69.180000  -8.145000  69.350000  -7.975000 ;
      RECT  69.250000 156.415000  69.420000 156.585000 ;
      RECT  69.540000  -8.145000  69.710000  -7.975000 ;
      RECT  69.610000 156.415000  69.780000 156.585000 ;
      RECT  69.900000  -8.145000  70.070000  -7.975000 ;
      RECT  69.970000 156.415000  70.140000 156.585000 ;
      RECT  70.260000  -8.145000  70.430000  -7.975000 ;
      RECT  70.330000 156.415000  70.500000 156.585000 ;
      RECT  70.620000  -8.145000  70.790000  -7.975000 ;
      RECT  70.690000 156.415000  70.860000 156.585000 ;
      RECT  70.980000  -8.145000  71.150000  -7.975000 ;
      RECT  71.050000 156.415000  71.220000 156.585000 ;
      RECT  71.340000  -8.145000  71.510000  -7.975000 ;
      RECT  71.410000 156.415000  71.580000 156.585000 ;
      RECT  71.700000  -8.145000  71.870000  -7.975000 ;
      RECT  71.770000 156.415000  71.940000 156.585000 ;
      RECT  72.060000  -8.145000  72.230000  -7.975000 ;
      RECT  72.130000 156.415000  72.300000 156.585000 ;
      RECT  72.420000  -8.145000  72.590000  -7.975000 ;
      RECT  72.490000 156.415000  72.660000 156.585000 ;
      RECT  72.780000  -8.145000  72.950000  -7.975000 ;
      RECT  72.850000 156.415000  73.020000 156.585000 ;
      RECT  73.140000  -8.145000  73.310000  -7.975000 ;
      RECT  73.210000 156.415000  73.380000 156.585000 ;
      RECT  73.500000  -8.145000  73.670000  -7.975000 ;
      RECT  73.570000 156.415000  73.740000 156.585000 ;
      RECT  73.860000  -8.145000  74.030000  -7.975000 ;
      RECT  73.930000 156.415000  74.100000 156.585000 ;
      RECT  74.220000  -8.145000  74.390000  -7.975000 ;
      RECT  74.290000 156.415000  74.460000 156.585000 ;
      RECT  74.580000  -8.145000  74.750000  -7.975000 ;
      RECT  74.650000 156.415000  74.820000 156.585000 ;
      RECT  74.940000  -8.145000  75.110000  -7.975000 ;
      RECT  75.010000 156.415000  75.180000 156.585000 ;
      RECT  75.300000  -8.145000  75.470000  -7.975000 ;
      RECT  75.370000 156.415000  75.540000 156.585000 ;
      RECT  75.660000  -8.145000  75.830000  -7.975000 ;
      RECT  75.730000 156.415000  75.900000 156.585000 ;
      RECT  76.020000  -8.145000  76.190000  -7.975000 ;
      RECT  76.090000 156.415000  76.260000 156.585000 ;
      RECT  76.380000  -8.145000  76.550000  -7.975000 ;
      RECT  76.450000 156.415000  76.620000 156.585000 ;
      RECT  76.740000  -8.145000  76.910000  -7.975000 ;
      RECT  76.810000 156.415000  76.980000 156.585000 ;
      RECT  77.100000  -8.145000  77.270000  -7.975000 ;
      RECT  77.175000 156.415000  77.345000 156.585000 ;
      RECT  77.460000  -8.145000  77.630000  -7.975000 ;
      RECT  77.540000 156.415000  77.710000 156.585000 ;
      RECT  77.820000  -8.145000  77.990000  -7.975000 ;
      RECT  77.905000 156.415000  78.075000 156.585000 ;
      RECT  78.180000  -8.145000  78.350000  -7.975000 ;
      RECT  78.270000 156.415000  78.440000 156.585000 ;
      RECT  78.540000  -8.145000  78.710000  -7.975000 ;
      RECT  78.635000 156.415000  78.805000 156.585000 ;
      RECT  78.900000  -8.145000  79.070000  -7.975000 ;
      RECT  79.000000 156.415000  79.170000 156.585000 ;
      RECT  79.260000  -8.145000  79.430000  -7.975000 ;
      RECT  79.365000 156.415000  79.535000 156.585000 ;
      RECT  79.620000  -8.145000  79.790000  -7.975000 ;
      RECT  79.730000 156.415000  79.900000 156.585000 ;
      RECT  79.980000  -8.145000  80.150000  -7.975000 ;
      RECT  80.095000 156.415000  80.265000 156.585000 ;
      RECT  80.340000  -8.145000  80.510000  -7.975000 ;
      RECT  80.460000 156.415000  80.630000 156.585000 ;
      RECT  80.700000  -8.145000  80.870000  -7.975000 ;
      RECT  80.825000 156.415000  80.995000 156.585000 ;
      RECT  81.060000  -8.145000  81.230000  -7.975000 ;
      RECT  81.190000 156.415000  81.360000 156.585000 ;
      RECT  81.420000  -8.145000  81.590000  -7.975000 ;
      RECT  81.555000 156.415000  81.725000 156.585000 ;
      RECT  81.780000  -8.145000  81.950000  -7.975000 ;
      RECT  81.920000 156.415000  82.090000 156.585000 ;
      RECT  82.140000  -8.145000  82.310000  -7.975000 ;
      RECT  82.285000 156.415000  82.455000 156.585000 ;
      RECT  82.500000  -8.145000  82.670000  -7.975000 ;
      RECT  82.650000 156.415000  82.820000 156.585000 ;
      RECT  82.860000  -8.145000  83.030000  -7.975000 ;
      RECT  83.015000 156.415000  83.185000 156.585000 ;
      RECT  83.220000  -8.145000  83.390000  -7.975000 ;
      RECT  83.380000 156.415000  83.550000 156.585000 ;
      RECT  83.580000  -8.145000  83.750000  -7.975000 ;
      RECT  83.745000 156.415000  83.915000 156.585000 ;
      RECT  83.940000  -8.145000  84.110000  -7.975000 ;
      RECT  84.110000 156.415000  84.280000 156.585000 ;
      RECT  84.300000  -8.145000  84.470000  -7.975000 ;
      RECT  84.475000 156.415000  84.645000 156.585000 ;
      RECT  84.660000  -8.145000  84.830000  -7.975000 ;
      RECT  84.840000 156.415000  85.010000 156.585000 ;
      RECT  85.020000  -8.145000  85.190000  -7.975000 ;
      RECT  85.205000 156.415000  85.375000 156.585000 ;
      RECT  85.380000  -8.145000  85.550000  -7.975000 ;
      RECT  85.570000 156.415000  85.740000 156.585000 ;
      RECT  85.740000  -8.145000  85.910000  -7.975000 ;
      RECT  85.935000 156.415000  86.105000 156.585000 ;
      RECT  86.100000  -8.145000  86.270000  -7.975000 ;
      RECT  86.300000 156.415000  86.470000 156.585000 ;
      RECT  86.460000  -8.145000  86.630000  -7.975000 ;
      RECT  86.665000 156.415000  86.835000 156.585000 ;
      RECT  86.820000  -8.145000  86.990000  -7.975000 ;
      RECT  87.030000 156.415000  87.200000 156.585000 ;
      RECT  87.180000  -8.145000  87.350000  -7.975000 ;
      RECT  87.395000 156.415000  87.565000 156.585000 ;
      RECT  87.540000  -8.145000  87.710000  -7.975000 ;
      RECT  87.760000 156.415000  87.930000 156.585000 ;
      RECT  87.900000  -8.145000  88.070000  -7.975000 ;
      RECT  88.125000 156.415000  88.295000 156.585000 ;
      RECT  88.260000  -8.145000  88.430000  -7.975000 ;
      RECT  88.490000 156.415000  88.660000 156.585000 ;
      RECT  88.620000  -8.145000  88.790000  -7.975000 ;
      RECT  88.855000 156.415000  89.025000 156.585000 ;
      RECT  88.980000  -8.145000  89.150000  -7.975000 ;
      RECT  89.220000 156.415000  89.390000 156.585000 ;
      RECT  89.340000  -8.145000  89.510000  -7.975000 ;
      RECT  89.585000 156.415000  89.755000 156.585000 ;
      RECT  89.700000  -8.145000  89.870000  -7.975000 ;
      RECT  89.950000 156.415000  90.120000 156.585000 ;
      RECT  90.060000  -8.145000  90.230000  -7.975000 ;
      RECT  90.315000 156.415000  90.485000 156.585000 ;
      RECT  90.420000  -8.145000  90.590000  -7.975000 ;
      RECT  90.680000 156.415000  90.850000 156.585000 ;
      RECT  90.780000  -8.145000  90.950000  -7.975000 ;
      RECT  91.045000 156.415000  91.215000 156.585000 ;
      RECT  91.140000  -8.145000  91.310000  -7.975000 ;
      RECT  91.410000 156.415000  91.580000 156.585000 ;
      RECT  91.500000  -8.145000  91.670000  -7.975000 ;
      RECT  91.775000 156.415000  91.945000 156.585000 ;
      RECT  91.860000  -8.145000  92.030000  -7.975000 ;
      RECT  92.140000 156.415000  92.310000 156.585000 ;
      RECT  92.220000  -8.145000  92.390000  -7.975000 ;
      RECT  92.505000 156.415000  92.675000 156.585000 ;
      RECT  92.580000  -8.145000  92.750000  -7.975000 ;
      RECT  92.870000 156.415000  93.040000 156.585000 ;
      RECT  92.940000  -8.145000  93.110000  -7.975000 ;
      RECT  93.235000 156.415000  93.405000 156.585000 ;
      RECT  93.300000  -8.145000  93.470000  -7.975000 ;
      RECT  93.600000 156.415000  93.770000 156.585000 ;
      RECT  93.660000  -8.145000  93.830000  -7.975000 ;
      RECT  93.965000 156.415000  94.135000 156.585000 ;
      RECT  94.020000  -8.145000  94.190000  -7.975000 ;
      RECT  94.330000 156.415000  94.500000 156.585000 ;
      RECT  94.380000  -8.145000  94.550000  -7.975000 ;
      RECT  94.695000 156.415000  94.865000 156.585000 ;
      RECT  94.740000  -8.145000  94.910000  -7.975000 ;
      RECT  95.060000 156.415000  95.230000 156.585000 ;
      RECT  95.100000  -8.145000  95.270000  -7.975000 ;
      RECT  95.425000 156.415000  95.595000 156.585000 ;
      RECT  95.460000  -8.145000  95.630000  -7.975000 ;
      RECT  95.790000 156.415000  95.960000 156.585000 ;
      RECT  95.820000  -8.145000  95.990000  -7.975000 ;
      RECT  96.155000 156.415000  96.325000 156.585000 ;
      RECT  96.180000  -8.145000  96.350000  -7.975000 ;
      RECT  96.520000 156.415000  96.690000 156.585000 ;
      RECT  96.540000  -8.145000  96.710000  -7.975000 ;
      RECT  96.885000 156.415000  97.055000 156.585000 ;
      RECT  96.900000  -8.145000  97.070000  -7.975000 ;
      RECT  97.250000 156.415000  97.420000 156.585000 ;
      RECT  97.260000  -8.145000  97.430000  -7.975000 ;
      RECT  97.615000 156.415000  97.785000 156.585000 ;
      RECT  97.620000  -8.145000  97.790000  -7.975000 ;
      RECT  97.980000 156.415000  98.150000 156.585000 ;
      RECT  98.065000  -8.060000  98.235000  -7.890000 ;
      RECT  98.065000  -7.695000  98.235000  -7.525000 ;
      RECT  98.065000  -7.330000  98.235000  -7.160000 ;
      RECT  98.065000  -6.965000  98.235000  -6.795000 ;
      RECT  98.065000  -6.600000  98.235000  -6.430000 ;
      RECT  98.065000  -6.235000  98.235000  -6.065000 ;
      RECT  98.065000  -5.870000  98.235000  -5.700000 ;
      RECT  98.065000  -5.505000  98.235000  -5.335000 ;
      RECT  98.065000  -5.140000  98.235000  -4.970000 ;
      RECT  98.065000  -4.775000  98.235000  -4.605000 ;
      RECT  98.065000  -4.410000  98.235000  -4.240000 ;
      RECT  98.065000  -4.045000  98.235000  -3.875000 ;
      RECT  98.065000  -3.680000  98.235000  -3.510000 ;
      RECT  98.065000  -3.315000  98.235000  -3.145000 ;
      RECT  98.065000  -2.950000  98.235000  -2.780000 ;
      RECT  98.065000  -2.585000  98.235000  -2.415000 ;
      RECT  98.065000  -2.220000  98.235000  -2.050000 ;
      RECT  98.065000  -1.855000  98.235000  -1.685000 ;
      RECT  98.065000  -1.490000  98.235000  -1.320000 ;
      RECT  98.065000  -1.125000  98.235000  -0.955000 ;
      RECT  98.065000  -0.760000  98.235000  -0.590000 ;
      RECT  98.065000  -0.395000  98.235000  -0.225000 ;
      RECT  98.065000  -0.030000  98.235000   0.140000 ;
      RECT  98.065000   0.335000  98.235000   0.505000 ;
      RECT  98.065000   0.700000  98.235000   0.870000 ;
      RECT  98.065000   1.065000  98.235000   1.235000 ;
      RECT  98.065000   1.430000  98.235000   1.600000 ;
      RECT  98.065000   1.795000  98.235000   1.965000 ;
      RECT  98.065000   2.160000  98.235000   2.330000 ;
      RECT  98.065000   2.525000  98.235000   2.695000 ;
      RECT  98.065000   2.890000  98.235000   3.060000 ;
      RECT  98.065000   3.255000  98.235000   3.425000 ;
      RECT  98.065000   3.620000  98.235000   3.790000 ;
      RECT  98.065000   3.985000  98.235000   4.155000 ;
      RECT  98.065000   4.350000  98.235000   4.520000 ;
      RECT  98.065000   4.715000  98.235000   4.885000 ;
      RECT  98.065000   5.080000  98.235000   5.250000 ;
      RECT  98.065000   5.445000  98.235000   5.615000 ;
      RECT  98.065000   5.810000  98.235000   5.980000 ;
      RECT  98.065000   6.175000  98.235000   6.345000 ;
      RECT  98.065000   6.540000  98.235000   6.710000 ;
      RECT  98.065000   6.905000  98.235000   7.075000 ;
      RECT  98.065000   7.270000  98.235000   7.440000 ;
      RECT  98.065000   7.635000  98.235000   7.805000 ;
      RECT  98.065000   8.000000  98.235000   8.170000 ;
      RECT  98.065000   8.365000  98.235000   8.535000 ;
      RECT  98.065000   8.730000  98.235000   8.900000 ;
      RECT  98.065000   9.090000  98.235000   9.260000 ;
      RECT  98.065000   9.450000  98.235000   9.620000 ;
      RECT  98.065000   9.810000  98.235000   9.980000 ;
      RECT  98.065000  10.170000  98.235000  10.340000 ;
      RECT  98.065000  10.530000  98.235000  10.700000 ;
      RECT  98.065000  10.890000  98.235000  11.060000 ;
      RECT  98.065000  11.250000  98.235000  11.420000 ;
      RECT  98.065000  11.610000  98.235000  11.780000 ;
      RECT  98.065000  11.970000  98.235000  12.140000 ;
      RECT  98.065000  12.330000  98.235000  12.500000 ;
      RECT  98.065000  12.690000  98.235000  12.860000 ;
      RECT  98.065000  13.050000  98.235000  13.220000 ;
      RECT  98.065000  13.410000  98.235000  13.580000 ;
      RECT  98.065000  13.770000  98.235000  13.940000 ;
      RECT  98.065000  14.130000  98.235000  14.300000 ;
      RECT  98.065000  14.490000  98.235000  14.660000 ;
      RECT  98.065000  14.850000  98.235000  15.020000 ;
      RECT  98.065000  15.210000  98.235000  15.380000 ;
      RECT  98.065000  15.570000  98.235000  15.740000 ;
      RECT  98.065000  15.930000  98.235000  16.100000 ;
      RECT  98.065000  16.290000  98.235000  16.460000 ;
      RECT  98.065000  16.650000  98.235000  16.820000 ;
      RECT  98.065000  17.010000  98.235000  17.180000 ;
      RECT  98.065000  17.370000  98.235000  17.540000 ;
      RECT  98.065000  17.730000  98.235000  17.900000 ;
      RECT  98.065000  18.090000  98.235000  18.260000 ;
      RECT  98.065000  18.450000  98.235000  18.620000 ;
      RECT  98.065000  18.810000  98.235000  18.980000 ;
      RECT  98.065000  19.170000  98.235000  19.340000 ;
      RECT  98.065000  19.530000  98.235000  19.700000 ;
      RECT  98.065000  19.890000  98.235000  20.060000 ;
      RECT  98.065000  20.250000  98.235000  20.420000 ;
      RECT  98.065000  20.610000  98.235000  20.780000 ;
      RECT  98.065000  20.970000  98.235000  21.140000 ;
      RECT  98.065000  21.330000  98.235000  21.500000 ;
      RECT  98.065000  21.690000  98.235000  21.860000 ;
      RECT  98.065000  22.050000  98.235000  22.220000 ;
      RECT  98.065000  22.410000  98.235000  22.580000 ;
      RECT  98.065000  22.770000  98.235000  22.940000 ;
      RECT  98.065000  23.130000  98.235000  23.300000 ;
      RECT  98.065000  23.490000  98.235000  23.660000 ;
      RECT  98.065000  23.850000  98.235000  24.020000 ;
      RECT  98.065000  24.210000  98.235000  24.380000 ;
      RECT  98.065000  24.570000  98.235000  24.740000 ;
      RECT  98.065000  24.930000  98.235000  25.100000 ;
      RECT  98.065000  25.290000  98.235000  25.460000 ;
      RECT  98.065000  25.650000  98.235000  25.820000 ;
      RECT  98.065000  26.010000  98.235000  26.180000 ;
      RECT  98.065000  26.370000  98.235000  26.540000 ;
      RECT  98.065000  26.730000  98.235000  26.900000 ;
      RECT  98.065000  27.090000  98.235000  27.260000 ;
      RECT  98.065000  27.450000  98.235000  27.620000 ;
      RECT  98.065000  27.810000  98.235000  27.980000 ;
      RECT  98.065000  28.170000  98.235000  28.340000 ;
      RECT  98.065000  28.530000  98.235000  28.700000 ;
      RECT  98.065000  28.890000  98.235000  29.060000 ;
      RECT  98.065000  29.250000  98.235000  29.420000 ;
      RECT  98.065000  29.610000  98.235000  29.780000 ;
      RECT  98.065000  29.970000  98.235000  30.140000 ;
      RECT  98.065000  30.330000  98.235000  30.500000 ;
      RECT  98.065000  30.690000  98.235000  30.860000 ;
      RECT  98.065000  31.050000  98.235000  31.220000 ;
      RECT  98.065000  31.410000  98.235000  31.580000 ;
      RECT  98.065000  31.770000  98.235000  31.940000 ;
      RECT  98.065000  32.130000  98.235000  32.300000 ;
      RECT  98.065000  32.490000  98.235000  32.660000 ;
      RECT  98.065000  32.850000  98.235000  33.020000 ;
      RECT  98.065000  33.210000  98.235000  33.380000 ;
      RECT  98.065000  33.570000  98.235000  33.740000 ;
      RECT  98.065000  33.930000  98.235000  34.100000 ;
      RECT  98.065000  34.290000  98.235000  34.460000 ;
      RECT  98.065000  34.650000  98.235000  34.820000 ;
      RECT  98.065000  35.010000  98.235000  35.180000 ;
      RECT  98.065000  35.370000  98.235000  35.540000 ;
      RECT  98.065000  35.730000  98.235000  35.900000 ;
      RECT  98.065000  36.090000  98.235000  36.260000 ;
      RECT  98.065000  36.450000  98.235000  36.620000 ;
      RECT  98.065000  36.810000  98.235000  36.980000 ;
      RECT  98.065000  37.170000  98.235000  37.340000 ;
      RECT  98.065000  37.530000  98.235000  37.700000 ;
      RECT  98.065000  37.890000  98.235000  38.060000 ;
      RECT  98.065000  38.250000  98.235000  38.420000 ;
      RECT  98.065000  38.610000  98.235000  38.780000 ;
      RECT  98.065000  38.970000  98.235000  39.140000 ;
      RECT  98.065000  39.330000  98.235000  39.500000 ;
      RECT  98.065000  39.690000  98.235000  39.860000 ;
      RECT  98.065000  40.050000  98.235000  40.220000 ;
      RECT  98.065000  40.410000  98.235000  40.580000 ;
      RECT  98.065000  40.770000  98.235000  40.940000 ;
      RECT  98.065000  41.130000  98.235000  41.300000 ;
      RECT  98.065000  41.490000  98.235000  41.660000 ;
      RECT  98.065000  41.850000  98.235000  42.020000 ;
      RECT  98.065000  42.210000  98.235000  42.380000 ;
      RECT  98.065000  42.570000  98.235000  42.740000 ;
      RECT  98.065000  42.930000  98.235000  43.100000 ;
      RECT  98.065000  43.290000  98.235000  43.460000 ;
      RECT  98.065000  43.650000  98.235000  43.820000 ;
      RECT  98.065000  44.010000  98.235000  44.180000 ;
      RECT  98.065000  44.370000  98.235000  44.540000 ;
      RECT  98.065000  44.730000  98.235000  44.900000 ;
      RECT  98.065000  45.090000  98.235000  45.260000 ;
      RECT  98.065000  45.450000  98.235000  45.620000 ;
      RECT  98.065000  45.810000  98.235000  45.980000 ;
      RECT  98.065000  46.170000  98.235000  46.340000 ;
      RECT  98.065000  46.530000  98.235000  46.700000 ;
      RECT  98.065000  46.890000  98.235000  47.060000 ;
      RECT  98.065000  47.250000  98.235000  47.420000 ;
      RECT  98.065000  47.610000  98.235000  47.780000 ;
      RECT  98.065000  47.970000  98.235000  48.140000 ;
      RECT  98.065000  48.330000  98.235000  48.500000 ;
      RECT  98.065000  48.690000  98.235000  48.860000 ;
      RECT  98.065000  49.050000  98.235000  49.220000 ;
      RECT  98.065000  49.410000  98.235000  49.580000 ;
      RECT  98.065000  49.770000  98.235000  49.940000 ;
      RECT  98.065000  50.130000  98.235000  50.300000 ;
      RECT  98.065000  50.490000  98.235000  50.660000 ;
      RECT  98.065000  50.850000  98.235000  51.020000 ;
      RECT  98.065000  51.210000  98.235000  51.380000 ;
      RECT  98.065000  51.570000  98.235000  51.740000 ;
      RECT  98.065000  51.930000  98.235000  52.100000 ;
      RECT  98.065000  52.290000  98.235000  52.460000 ;
      RECT  98.065000  52.650000  98.235000  52.820000 ;
      RECT  98.065000  53.010000  98.235000  53.180000 ;
      RECT  98.065000  53.370000  98.235000  53.540000 ;
      RECT  98.065000  53.730000  98.235000  53.900000 ;
      RECT  98.065000  54.090000  98.235000  54.260000 ;
      RECT  98.065000  54.450000  98.235000  54.620000 ;
      RECT  98.065000  54.810000  98.235000  54.980000 ;
      RECT  98.065000  55.170000  98.235000  55.340000 ;
      RECT  98.065000  55.530000  98.235000  55.700000 ;
      RECT  98.065000  55.890000  98.235000  56.060000 ;
      RECT  98.065000  56.250000  98.235000  56.420000 ;
      RECT  98.065000  56.610000  98.235000  56.780000 ;
      RECT  98.065000  56.970000  98.235000  57.140000 ;
      RECT  98.065000  57.330000  98.235000  57.500000 ;
      RECT  98.065000  57.690000  98.235000  57.860000 ;
      RECT  98.065000  58.050000  98.235000  58.220000 ;
      RECT  98.065000  58.410000  98.235000  58.580000 ;
      RECT  98.065000  58.770000  98.235000  58.940000 ;
      RECT  98.065000  59.130000  98.235000  59.300000 ;
      RECT  98.065000  59.490000  98.235000  59.660000 ;
      RECT  98.065000  59.850000  98.235000  60.020000 ;
      RECT  98.065000  60.210000  98.235000  60.380000 ;
      RECT  98.065000  60.570000  98.235000  60.740000 ;
      RECT  98.065000  60.930000  98.235000  61.100000 ;
      RECT  98.065000  61.290000  98.235000  61.460000 ;
      RECT  98.065000  61.650000  98.235000  61.820000 ;
      RECT  98.065000  62.010000  98.235000  62.180000 ;
      RECT  98.065000  62.370000  98.235000  62.540000 ;
      RECT  98.065000  62.730000  98.235000  62.900000 ;
      RECT  98.065000  63.090000  98.235000  63.260000 ;
      RECT  98.065000  63.450000  98.235000  63.620000 ;
      RECT  98.065000  63.810000  98.235000  63.980000 ;
      RECT  98.065000  64.170000  98.235000  64.340000 ;
      RECT  98.065000  64.530000  98.235000  64.700000 ;
      RECT  98.065000  64.890000  98.235000  65.060000 ;
      RECT  98.065000  65.250000  98.235000  65.420000 ;
      RECT  98.065000  65.610000  98.235000  65.780000 ;
      RECT  98.065000  65.970000  98.235000  66.140000 ;
      RECT  98.065000  66.330000  98.235000  66.500000 ;
      RECT  98.065000  66.690000  98.235000  66.860000 ;
      RECT  98.065000  67.050000  98.235000  67.220000 ;
      RECT  98.065000  67.410000  98.235000  67.580000 ;
      RECT  98.065000  67.770000  98.235000  67.940000 ;
      RECT  98.065000  68.130000  98.235000  68.300000 ;
      RECT  98.065000  68.490000  98.235000  68.660000 ;
      RECT  98.065000  68.850000  98.235000  69.020000 ;
      RECT  98.065000  69.210000  98.235000  69.380000 ;
      RECT  98.065000  69.570000  98.235000  69.740000 ;
      RECT  98.065000  69.930000  98.235000  70.100000 ;
      RECT  98.065000  70.290000  98.235000  70.460000 ;
      RECT  98.065000  70.650000  98.235000  70.820000 ;
      RECT  98.065000  71.010000  98.235000  71.180000 ;
      RECT  98.065000  71.370000  98.235000  71.540000 ;
      RECT  98.065000  71.730000  98.235000  71.900000 ;
      RECT  98.065000  72.090000  98.235000  72.260000 ;
      RECT  98.065000  72.450000  98.235000  72.620000 ;
      RECT  98.065000  72.810000  98.235000  72.980000 ;
      RECT  98.065000  73.170000  98.235000  73.340000 ;
      RECT  98.065000  73.530000  98.235000  73.700000 ;
      RECT  98.065000  73.890000  98.235000  74.060000 ;
      RECT  98.065000  74.250000  98.235000  74.420000 ;
      RECT  98.065000  74.610000  98.235000  74.780000 ;
      RECT  98.065000  74.970000  98.235000  75.140000 ;
      RECT  98.065000  75.330000  98.235000  75.500000 ;
      RECT  98.065000  75.690000  98.235000  75.860000 ;
      RECT  98.065000  76.050000  98.235000  76.220000 ;
      RECT  98.065000  76.410000  98.235000  76.580000 ;
      RECT  98.065000  76.770000  98.235000  76.940000 ;
      RECT  98.065000  77.130000  98.235000  77.300000 ;
      RECT  98.065000  77.490000  98.235000  77.660000 ;
      RECT  98.065000  77.850000  98.235000  78.020000 ;
      RECT  98.065000  78.210000  98.235000  78.380000 ;
      RECT  98.065000  78.570000  98.235000  78.740000 ;
      RECT  98.065000  78.930000  98.235000  79.100000 ;
      RECT  98.065000  79.290000  98.235000  79.460000 ;
      RECT  98.065000  79.650000  98.235000  79.820000 ;
      RECT  98.065000  80.010000  98.235000  80.180000 ;
      RECT  98.065000  80.370000  98.235000  80.540000 ;
      RECT  98.065000  80.730000  98.235000  80.900000 ;
      RECT  98.065000  81.090000  98.235000  81.260000 ;
      RECT  98.065000  81.450000  98.235000  81.620000 ;
      RECT  98.065000  81.810000  98.235000  81.980000 ;
      RECT  98.065000  82.170000  98.235000  82.340000 ;
      RECT  98.065000  82.530000  98.235000  82.700000 ;
      RECT  98.065000  82.890000  98.235000  83.060000 ;
      RECT  98.065000  83.250000  98.235000  83.420000 ;
      RECT  98.065000  83.610000  98.235000  83.780000 ;
      RECT  98.065000  83.970000  98.235000  84.140000 ;
      RECT  98.065000  84.330000  98.235000  84.500000 ;
      RECT  98.065000  84.690000  98.235000  84.860000 ;
      RECT  98.065000  85.050000  98.235000  85.220000 ;
      RECT  98.065000  85.410000  98.235000  85.580000 ;
      RECT  98.065000  85.770000  98.235000  85.940000 ;
      RECT  98.065000  86.130000  98.235000  86.300000 ;
      RECT  98.065000  86.490000  98.235000  86.660000 ;
      RECT  98.065000  86.850000  98.235000  87.020000 ;
      RECT  98.065000  87.210000  98.235000  87.380000 ;
      RECT  98.065000  87.570000  98.235000  87.740000 ;
      RECT  98.065000  87.930000  98.235000  88.100000 ;
      RECT  98.065000  88.290000  98.235000  88.460000 ;
      RECT  98.065000  88.650000  98.235000  88.820000 ;
      RECT  98.065000  89.010000  98.235000  89.180000 ;
      RECT  98.065000  89.370000  98.235000  89.540000 ;
      RECT  98.065000  89.730000  98.235000  89.900000 ;
      RECT  98.065000  90.090000  98.235000  90.260000 ;
      RECT  98.065000  90.450000  98.235000  90.620000 ;
      RECT  98.065000  90.810000  98.235000  90.980000 ;
      RECT  98.065000  91.170000  98.235000  91.340000 ;
      RECT  98.065000  91.530000  98.235000  91.700000 ;
      RECT  98.065000  91.890000  98.235000  92.060000 ;
      RECT  98.065000  92.250000  98.235000  92.420000 ;
      RECT  98.065000  92.610000  98.235000  92.780000 ;
      RECT  98.065000  92.970000  98.235000  93.140000 ;
      RECT  98.065000  93.330000  98.235000  93.500000 ;
      RECT  98.065000  93.690000  98.235000  93.860000 ;
      RECT  98.065000  94.050000  98.235000  94.220000 ;
      RECT  98.065000  94.410000  98.235000  94.580000 ;
      RECT  98.065000  94.770000  98.235000  94.940000 ;
      RECT  98.065000  95.130000  98.235000  95.300000 ;
      RECT  98.065000  95.490000  98.235000  95.660000 ;
      RECT  98.065000  95.850000  98.235000  96.020000 ;
      RECT  98.065000  96.210000  98.235000  96.380000 ;
      RECT  98.065000  96.570000  98.235000  96.740000 ;
      RECT  98.065000  96.930000  98.235000  97.100000 ;
      RECT  98.065000  97.290000  98.235000  97.460000 ;
      RECT  98.065000  97.650000  98.235000  97.820000 ;
      RECT  98.065000  98.010000  98.235000  98.180000 ;
      RECT  98.065000  98.370000  98.235000  98.540000 ;
      RECT  98.065000  98.730000  98.235000  98.900000 ;
      RECT  98.065000  99.090000  98.235000  99.260000 ;
      RECT  98.065000  99.450000  98.235000  99.620000 ;
      RECT  98.065000  99.810000  98.235000  99.980000 ;
      RECT  98.065000 100.170000  98.235000 100.340000 ;
      RECT  98.065000 100.530000  98.235000 100.700000 ;
      RECT  98.065000 100.890000  98.235000 101.060000 ;
      RECT  98.065000 101.250000  98.235000 101.420000 ;
      RECT  98.065000 101.610000  98.235000 101.780000 ;
      RECT  98.065000 101.970000  98.235000 102.140000 ;
      RECT  98.065000 102.330000  98.235000 102.500000 ;
      RECT  98.065000 102.690000  98.235000 102.860000 ;
      RECT  98.065000 103.050000  98.235000 103.220000 ;
      RECT  98.065000 103.410000  98.235000 103.580000 ;
      RECT  98.065000 103.770000  98.235000 103.940000 ;
      RECT  98.065000 104.130000  98.235000 104.300000 ;
      RECT  98.065000 104.490000  98.235000 104.660000 ;
      RECT  98.065000 104.850000  98.235000 105.020000 ;
      RECT  98.065000 105.210000  98.235000 105.380000 ;
      RECT  98.065000 105.570000  98.235000 105.740000 ;
      RECT  98.065000 105.930000  98.235000 106.100000 ;
      RECT  98.065000 106.290000  98.235000 106.460000 ;
      RECT  98.065000 106.650000  98.235000 106.820000 ;
      RECT  98.065000 107.010000  98.235000 107.180000 ;
      RECT  98.065000 107.370000  98.235000 107.540000 ;
      RECT  98.065000 107.730000  98.235000 107.900000 ;
      RECT  98.065000 108.090000  98.235000 108.260000 ;
      RECT  98.065000 108.450000  98.235000 108.620000 ;
      RECT  98.065000 108.810000  98.235000 108.980000 ;
      RECT  98.065000 109.170000  98.235000 109.340000 ;
      RECT  98.065000 109.530000  98.235000 109.700000 ;
      RECT  98.065000 109.890000  98.235000 110.060000 ;
      RECT  98.065000 110.250000  98.235000 110.420000 ;
      RECT  98.065000 110.610000  98.235000 110.780000 ;
      RECT  98.065000 110.970000  98.235000 111.140000 ;
      RECT  98.065000 111.330000  98.235000 111.500000 ;
      RECT  98.065000 111.690000  98.235000 111.860000 ;
      RECT  98.065000 112.050000  98.235000 112.220000 ;
      RECT  98.065000 112.410000  98.235000 112.580000 ;
      RECT  98.065000 112.770000  98.235000 112.940000 ;
      RECT  98.065000 113.130000  98.235000 113.300000 ;
      RECT  98.065000 113.490000  98.235000 113.660000 ;
      RECT  98.065000 113.850000  98.235000 114.020000 ;
      RECT  98.065000 114.210000  98.235000 114.380000 ;
      RECT  98.065000 114.570000  98.235000 114.740000 ;
      RECT  98.065000 114.930000  98.235000 115.100000 ;
      RECT  98.065000 115.290000  98.235000 115.460000 ;
      RECT  98.065000 115.650000  98.235000 115.820000 ;
      RECT  98.065000 116.010000  98.235000 116.180000 ;
      RECT  98.065000 116.370000  98.235000 116.540000 ;
      RECT  98.065000 116.730000  98.235000 116.900000 ;
      RECT  98.065000 117.090000  98.235000 117.260000 ;
      RECT  98.065000 117.450000  98.235000 117.620000 ;
      RECT  98.065000 117.810000  98.235000 117.980000 ;
      RECT  98.065000 118.170000  98.235000 118.340000 ;
      RECT  98.065000 118.530000  98.235000 118.700000 ;
      RECT  98.065000 118.890000  98.235000 119.060000 ;
      RECT  98.065000 119.250000  98.235000 119.420000 ;
      RECT  98.065000 119.610000  98.235000 119.780000 ;
      RECT  98.065000 119.970000  98.235000 120.140000 ;
      RECT  98.065000 120.330000  98.235000 120.500000 ;
      RECT  98.065000 120.690000  98.235000 120.860000 ;
      RECT  98.065000 121.050000  98.235000 121.220000 ;
      RECT  98.065000 121.410000  98.235000 121.580000 ;
      RECT  98.065000 121.770000  98.235000 121.940000 ;
      RECT  98.065000 122.130000  98.235000 122.300000 ;
      RECT  98.065000 122.490000  98.235000 122.660000 ;
      RECT  98.065000 122.850000  98.235000 123.020000 ;
      RECT  98.065000 123.210000  98.235000 123.380000 ;
      RECT  98.065000 123.570000  98.235000 123.740000 ;
      RECT  98.065000 123.930000  98.235000 124.100000 ;
      RECT  98.065000 124.290000  98.235000 124.460000 ;
      RECT  98.065000 124.650000  98.235000 124.820000 ;
      RECT  98.065000 125.010000  98.235000 125.180000 ;
      RECT  98.065000 125.370000  98.235000 125.540000 ;
      RECT  98.065000 125.730000  98.235000 125.900000 ;
      RECT  98.065000 126.090000  98.235000 126.260000 ;
      RECT  98.065000 126.450000  98.235000 126.620000 ;
      RECT  98.065000 126.810000  98.235000 126.980000 ;
      RECT  98.065000 127.170000  98.235000 127.340000 ;
      RECT  98.065000 127.530000  98.235000 127.700000 ;
      RECT  98.065000 127.890000  98.235000 128.060000 ;
      RECT  98.065000 128.250000  98.235000 128.420000 ;
      RECT  98.065000 128.610000  98.235000 128.780000 ;
      RECT  98.065000 128.970000  98.235000 129.140000 ;
      RECT  98.065000 129.330000  98.235000 129.500000 ;
      RECT  98.065000 129.690000  98.235000 129.860000 ;
      RECT  98.065000 130.050000  98.235000 130.220000 ;
      RECT  98.065000 130.410000  98.235000 130.580000 ;
      RECT  98.065000 130.770000  98.235000 130.940000 ;
      RECT  98.065000 131.130000  98.235000 131.300000 ;
      RECT  98.065000 131.490000  98.235000 131.660000 ;
      RECT  98.065000 131.850000  98.235000 132.020000 ;
      RECT  98.065000 132.210000  98.235000 132.380000 ;
      RECT  98.065000 132.570000  98.235000 132.740000 ;
      RECT  98.065000 132.930000  98.235000 133.100000 ;
      RECT  98.065000 133.290000  98.235000 133.460000 ;
      RECT  98.065000 133.650000  98.235000 133.820000 ;
      RECT  98.065000 134.010000  98.235000 134.180000 ;
      RECT  98.065000 134.370000  98.235000 134.540000 ;
      RECT  98.065000 134.730000  98.235000 134.900000 ;
      RECT  98.065000 135.090000  98.235000 135.260000 ;
      RECT  98.065000 135.450000  98.235000 135.620000 ;
      RECT  98.065000 135.810000  98.235000 135.980000 ;
      RECT  98.065000 136.170000  98.235000 136.340000 ;
      RECT  98.065000 136.530000  98.235000 136.700000 ;
      RECT  98.065000 136.890000  98.235000 137.060000 ;
      RECT  98.065000 137.250000  98.235000 137.420000 ;
      RECT  98.065000 137.610000  98.235000 137.780000 ;
      RECT  98.065000 137.970000  98.235000 138.140000 ;
      RECT  98.065000 138.330000  98.235000 138.500000 ;
      RECT  98.065000 138.690000  98.235000 138.860000 ;
      RECT  98.065000 139.050000  98.235000 139.220000 ;
      RECT  98.065000 139.410000  98.235000 139.580000 ;
      RECT  98.065000 139.770000  98.235000 139.940000 ;
      RECT  98.065000 140.130000  98.235000 140.300000 ;
      RECT  98.065000 140.490000  98.235000 140.660000 ;
      RECT  98.065000 140.850000  98.235000 141.020000 ;
      RECT  98.065000 141.210000  98.235000 141.380000 ;
      RECT  98.065000 141.570000  98.235000 141.740000 ;
      RECT  98.065000 141.930000  98.235000 142.100000 ;
      RECT  98.065000 142.290000  98.235000 142.460000 ;
      RECT  98.065000 142.650000  98.235000 142.820000 ;
      RECT  98.065000 143.010000  98.235000 143.180000 ;
      RECT  98.065000 143.370000  98.235000 143.540000 ;
      RECT  98.065000 143.730000  98.235000 143.900000 ;
      RECT  98.065000 144.090000  98.235000 144.260000 ;
      RECT  98.065000 144.450000  98.235000 144.620000 ;
      RECT  98.065000 144.810000  98.235000 144.980000 ;
      RECT  98.065000 145.170000  98.235000 145.340000 ;
      RECT  98.065000 145.530000  98.235000 145.700000 ;
      RECT  98.065000 145.890000  98.235000 146.060000 ;
      RECT  98.065000 146.250000  98.235000 146.420000 ;
      RECT  98.065000 146.610000  98.235000 146.780000 ;
      RECT  98.065000 146.970000  98.235000 147.140000 ;
      RECT  98.065000 147.330000  98.235000 147.500000 ;
      RECT  98.065000 147.690000  98.235000 147.860000 ;
      RECT  98.065000 148.050000  98.235000 148.220000 ;
      RECT  98.065000 148.410000  98.235000 148.580000 ;
      RECT  98.065000 148.770000  98.235000 148.940000 ;
      RECT  98.065000 149.130000  98.235000 149.300000 ;
      RECT  98.065000 149.490000  98.235000 149.660000 ;
      RECT  98.065000 149.850000  98.235000 150.020000 ;
      RECT  98.065000 150.210000  98.235000 150.380000 ;
      RECT  98.065000 150.570000  98.235000 150.740000 ;
      RECT  98.065000 150.930000  98.235000 151.100000 ;
      RECT  98.065000 151.290000  98.235000 151.460000 ;
      RECT  98.065000 151.650000  98.235000 151.820000 ;
      RECT  98.065000 152.010000  98.235000 152.180000 ;
      RECT  98.065000 152.370000  98.235000 152.540000 ;
      RECT  98.065000 152.730000  98.235000 152.900000 ;
      RECT  98.065000 153.090000  98.235000 153.260000 ;
      RECT  98.065000 153.450000  98.235000 153.620000 ;
      RECT  98.065000 153.810000  98.235000 153.980000 ;
      RECT  98.065000 154.170000  98.235000 154.340000 ;
      RECT  98.065000 154.530000  98.235000 154.700000 ;
      RECT  98.065000 154.890000  98.235000 155.060000 ;
      RECT  98.065000 155.250000  98.235000 155.420000 ;
      RECT  98.065000 155.610000  98.235000 155.780000 ;
      RECT  98.065000 155.970000  98.235000 156.140000 ;
    LAYER met1 ;
      RECT -98.300000  -8.210000  98.300000  -7.910000 ;
      RECT -98.300000  -7.910000 -98.000000 156.350000 ;
      RECT -98.300000 156.350000  98.300000 156.650000 ;
      RECT  -2.700000  -6.910000   2.700000 155.350000 ;
      RECT  98.000000  -7.910000  98.300000 156.350000 ;
    LAYER met2 ;
      RECT -1.985000 2.960000 1.985000 4.490000 ;
    LAYER met3 ;
      RECT -2.000000 2.870000 2.000000 47.495000 ;
    LAYER met4 ;
      POLYGON  -5.240000  17.495000 -2.760000  17.495000 -2.760000  15.015000 ;
      POLYGON  -5.240000  33.495000 -2.760000  33.495000 -2.760000  31.015000 ;
      POLYGON  -3.240000 108.495000 -3.240000 106.495000 -5.240000 106.495000 ;
      POLYGON  -3.240000 124.495000 -3.240000 122.495000 -5.240000 122.495000 ;
      POLYGON  -3.240000 140.495000 -3.240000 138.495000 -5.240000 138.495000 ;
      POLYGON  -2.760000  15.015000  2.760000  15.015000  2.760000   9.495000 ;
      POLYGON  -2.760000  23.495000  5.240000  15.495000 -2.760000  15.495000 ;
      POLYGON  -2.760000  31.015000  2.760000  31.015000  2.760000  25.495000 ;
      POLYGON  -2.760000  39.495000  5.240000  31.495000 -2.760000  31.495000 ;
      POLYGON  -2.760000 108.495000  5.240000 108.495000 -2.760000 100.495000 ;
      POLYGON  -2.760000 124.495000  5.240000 124.495000 -2.760000 116.495000 ;
      POLYGON  -2.760000 140.495000  5.240000 140.495000 -2.760000 132.495000 ;
      POLYGON   2.760000 114.495000  2.760000 108.495000 -3.240000 108.495000 ;
      POLYGON   2.760000 130.495000  2.760000 124.495000 -3.240000 124.495000 ;
      POLYGON   2.760000 146.495000  2.760000 140.495000 -3.240000 140.495000 ;
      RECT -16.080000  17.495000 -2.760000  23.495000 ;
      RECT -16.080000  33.495000 -2.760000  39.495000 ;
      RECT -16.080000 100.495000 -2.760000 106.495000 ;
      RECT -16.080000 116.495000 -2.760000 122.495000 ;
      RECT -16.080000 132.495000 -2.760000 138.495000 ;
      RECT  -3.240000 106.495000 -2.760000 108.495000 ;
      RECT  -3.240000 122.495000 -2.760000 124.495000 ;
      RECT  -3.240000 138.495000 -2.760000 140.495000 ;
      RECT  -2.760000  15.015000 16.080000  15.495000 ;
      RECT  -2.760000  31.015000 16.080000  31.495000 ;
      RECT  -1.795000  41.910000  1.785000  47.040000 ;
      RECT   2.760000   9.495000 16.080000  15.015000 ;
      RECT   2.760000  25.495000 16.080000  31.015000 ;
      RECT   2.760000 108.495000 16.080000 114.495000 ;
      RECT   2.760000 124.495000 16.080000 130.495000 ;
      RECT   2.760000 140.495000 16.080000 146.495000 ;
    LAYER via2 ;
      RECT -1.940000 2.985000 1.940000 4.465000 ;
    LAYER via3 ;
      RECT -1.765000 41.915000 1.755000 47.035000 ;
    LAYER via4 ;
      RECT -15.670000  18.305000 -6.490000  22.685000 ;
      RECT -15.670000  34.305000 -6.490000  38.685000 ;
      RECT -15.670000 101.305000 -6.490000 105.685000 ;
      RECT -15.670000 117.305000 -6.490000 121.685000 ;
      RECT -15.670000 133.305000 -6.490000 137.685000 ;
      RECT  -1.420000  42.285000  1.360000  46.665000 ;
      RECT   6.490000  10.305000 15.670000  14.685000 ;
      RECT   6.490000  26.305000 15.670000  30.685000 ;
      RECT   6.490000 109.305000 15.670000 113.685000 ;
      RECT   6.490000 125.305000 15.670000 129.685000 ;
      RECT   6.490000 141.305000 15.670000 145.685000 ;
  END
END sky130_fd_pr__ind_01_04
END LIBRARY
