* SKY130 legacy discrete models
* Parameters used by res_generic_nd/pd__hv
.param
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = 9.3222e-1
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = 9.4436e-1
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = 1.1726e+0
+ sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult = 1.2510e+0

.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_nfet_01v8__fs.corner.spice"
