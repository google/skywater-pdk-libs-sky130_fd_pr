# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__res_high_po_1p41__example1
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__res_high_po_1p41__example1 ;
  ORIGIN  2.080000  0.000000 ;
  SIZE  5.570000 BY  1.410000 ;
  OBS
    LAYER li1 ;
      RECT -2.080000 0.000000 0.060000 0.180000 ;
      RECT -2.080000 0.180000 0.080000 1.230000 ;
      RECT -2.080000 1.230000 0.060000 1.410000 ;
      RECT  1.330000 0.180000 3.490000 1.230000 ;
      RECT  1.350000 0.000000 3.490000 0.180000 ;
      RECT  1.350000 1.230000 3.490000 1.410000 ;
    LAYER mcon ;
      RECT -1.970000 0.260000 0.000000 1.150000 ;
      RECT  1.410000 0.260000 3.380000 1.150000 ;
    LAYER met1 ;
      RECT -2.030000 0.200000 0.060000 1.210000 ;
      RECT  1.350000 0.200000 3.440000 1.210000 ;
  END
END sky130_fd_pr__res_high_po_1p41__example1
END LIBRARY
