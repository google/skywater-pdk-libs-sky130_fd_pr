* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* ./models_bjt.spice created from ./models.spice
*
**********************************
******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/04/05  UZMN (Usman Suriono)
*      Why     : New infrastructure of an npn model
*      What    : Converted from  nsky130_fd_pr__pnp_05v5_W0p68L0p68ar1x1 model
*                Replaced all junction capacitance variation by correlated diodes.

.subckt  sky130_fd_pr__npn_05v5_W1p00L1p00 c b e s mult=1
+
+ 
.param  dkisnpn1x1 = 8.7913e-01
+ dkbfnpn1x1 = 9.8501e-01
+ var_is = {1/sw_func_rdn**2*(1+1.58*sw_mm_npn_is*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}
+ var_bf = {(sw_func_pw_rs*sw_pw_rs_mc)**2.2*(1+1.05*sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}


Qsky130_fd_pr__npn_05v5_W1p00L1p00 c b e s sky130_fd_pr__npn_05v5_W1p00L1p00_model 



.model sky130_fd_pr__npn_05v5_W1p00L1p00_model npn level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ dcap = 2
+ cjc = '1.73302e-014*sw_func_pw_dnw_cj'
+ cje = '5.4899e-015*sw_func_nsd_pw_cj'
+ cjs = '3.03477e-014*sw_func_dnw_sub_cj'
+ fc = 0.5 mjc = 0.33982 mje = 0.44
+ mjs = 0.49 vjc = 0.58758 vje = 0.729 vjs = 0.5348
+ xcjc = 1 itf = '2.6e-03+4e-3' ptf = 20 tf = '7.24041e-011+2e-11'
+ tr = 0 vtf = '0.5+0.2' xtf = '2.0-0.9'
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.523963 kf = 6.1811298e-11
**************************************************************
*               DC PARAMETERS
**************************************************************
+ is = '4.5584e-018*dkisnpn1x1*var_is'
+ bf = '39.28*dkbfnpn1x1*var_bf'
+ ise = '3.2947e-016*(1-sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))'
+ vaf = '100 / var_bf'
+ subs = 1 rb = 602.54 re = 30
+ irb = 7.4e+020 rc = 320.4 rbm = 0
+ nf = 1.0394 ikf = 0.00083757
+ ne = 1.792 ns = 1.0 br = 1 ibc = 0
+ iss = 0 nr = 0.8976 var = 0 ikr = 3.679e-07
+ nkf = 0.5 isc = 0 nc = 2
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xtb = 0 xti = 1.0713 eg = 1.188 gap1 = 0
+ gap2 = 0 ctc = 0
+ cte = 0 cts = 0 tlev = 0 tlevc = 0
+ tvjc = 0 tvje = 0 tvjs = 0
+ tis1 = 0 tise1 = 0 tisc1 = 0
+ tnf1 = 4.208e-005 tnr1 = -0.0011234 tne1 = 0 tnc1 = 0
+ tbf1 = 0.00776 tbr1 = 0 tiss1 = 0 tvaf1 = 0
+ tvar1 = 0 tikf1 = -0.0074 tikr1 = 0 tns1 = 0
+ trb1 = 0 trc1 = 0 tre1 = 0 tirb1 = 0
+ tsky130_fd_pr__res_generic_m1 = 0 tmjc1 = 0 tmje1 = 0 tmjs1 = 0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 4e-012
+ tise2 = 0 tisc2 = 0 tnf2 = -3.372e-007
+ tnr2 = -2.274e-006
+ tne2 = 0 tnc2 = 0 tbf2 = 6.48e-006 tbr2 = 0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 4e-005
+ tikr2 = 0 tns2 = 0 trb2 = 0 trc2 = 0
+ tre2 = 0 tirb2 = 0 tsky130_fd_pr__res_generic_m2 = 0 tmjc2 = 0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0
**************************************************************
*               QUASI
**************************************************************

.ends sky130_fd_pr__npn_05v5_W1p00L1p00

******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/02/20  UZMN (Usman Suriono)
*      Why     : New infrastructure of an npn model
*      What    : Converted from  sky130_fd_pr__npn_05v5_W1p00L1p00_2p0_hv model
*                Replaced all junction capacitance variation by correlated diodes.


.subckt  sky130_fd_pr__npn_11v0_W1p00L1p00 c b e s mult=1

+
+ 
.param  var_is = {1/sw_func_rdn**2*(1+sw_mm_npn_is*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}
+ var_bf = {(sw_func_pw_rs*sw_pw_rs_mc)**2.6*(1+sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}

rc c c1 r = 440 tc1 = -4e-3
q2 s c1 b s sky130_fd_pr__pnp_05v5_W0p68L0p68_polyhv 
xd1 s b sky130_fd_pr__model__parasitic__diode_ps2dn area = 1.34 perim = 0.6
Qsky130_fd_pr__npn_11v0_W1p00L1p00 c1 b e s sky130_fd_pr__npn_11v0_W1p00L1p00_base 


.model sky130_fd_pr__npn_11v0_W1p00L1p00_base npn level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ dcap = 2
+ cjc = '1.60339e-014*sw_func_pw_dnw_cj'
+ cje = '10.30981e-015*sw_func_nsd_pw_cj'
+ cjs = '3.05951e-014*sw_func_dnw_sub_cj'
+ fc = 0.5 mjc = 0.33982 mje = 0.44
+ mjs = 0.49 vjc = 0.58758 vje = 0.729 vjs = 0.5348
+ xcjc = 1 itf = 9.6e-03 ptf = 20 tf = 10.84e-011
+ tr = 0 vtf = 0.5 xtf = 2.9
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.9 kf = 5.0e-010
**************************************************************
*               DC PARAMETERS
**************************************************************
+ is = '1.1082e-017*var_is'
+ bf = '141.286*var_bf'
+ ise = '5.3935e-016*(1-sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))'
+ vaf = '100 / var_bf'
+ ikf = 0.00046731
+ nf = 1.0262306
+ rb = 1400
+ re = 85 irb = 4.424e-005 rc = 1.0 rbm = 400.07
+ ne = 1.7527 ns = 1 br = 100
+ iss = 0 nr = 1.0262306
+ var = 0 ikr = 0.00046731 nkf = 0.31875 isc = 0
+ nc = 2
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xtb = 0 xti = 2.7498 eg = 1.1714 gap1 = 0
+ gap2 = 0 ctc = 0 cte = 0 cts = 0
+ tlev = 0 tlevc = 0 tvjc = 0 tvje = 0
+ tvjs = 0 tis1 = 0 tise1 = 0 tisc1 = 0
+ tnf1 = 4.208e-005 tnr1 = -0.000522 tne1 = 0 tnc1 = 0
+ tbf1 = 7.4942e-003 tbr1 = 0 tiss1 = 0 tvaf1 = 0
+ tvar1 = 0 tikf1 = -0.012219846 tikr1 = 0 tns1 = 0
+ trb1 = -0.0029419354 trc1 = 3.7260032e-005 tre1 = 5e-3 tirb1 = 0
+ tsky130_fd_pr__res_generic_m1 = 0.004459028 tmjc1 = 0 tmje1 = 0 tmjs1 = 0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 4e-012
+ tise2 = 0 tisc2 = 0 tnf2 = -3.372e-007 tnr2 = 1.8e-006
+ tne2 = 0 tnc2 = 0 tbf2 = 7.633e-006 tbr2 = 0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 9.3646292e-005
+ tikr2 = 0 tns2 = 0 trb2 = 3.4143764e-005 trc2 = 3.0650517e-007
+ tre2 = 0.0 tirb2 = 0 tsky130_fd_pr__res_generic_m2 = -4.9458296e-005 tmjc2 = 0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0 titf2 = 0
+ ttr2 = 0
**************************************************************
*               QUASI
**************************************************************
**


.model sky130_fd_pr__pnp_05v5_W0p68L0p68_polyhv pnp level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ dcap = 2 cjc = 0 cje = 0
+ cjs = 0 fc = 0.5 mjc = 0.33 mje = 0.33
+ mjs = 0.5 vjc = 0.75 vje = 0.75 vjs = 0.75
+ xcjc = 1
+ itf = 0 ptf = 0 tf = 0 tr = 0
+ vtf = 0.5 xtf = 0
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.9 kf = 5.0e-09
**************************************************************
*               DC PARAMETERS
**************************************************************
+ is = '1.2252871e-016*var_is'
+ bf = '25*var_bf'
+ nf = 1.0161516 vaf = 0 ikf = 100
+ rb = 1922.4
+ re = 6000 irb = 0 rc = 1 rbm = 46.144
+ ise = 1e-016 ne = 2 ns = 1 br = 1
+ ibc = 0 iss = 0 nr = 1
+ var = 0 ikr = 1e-10 nkf = 0.41826 isc = 0
+ nc = 2
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xtb = 0 xti = 5.351377 eg = 1.11 gap1 = 0
+ gap2 = 0 ctc = 0
+ cte = 0 cts = 0 tlev = 0 tlevc = 0
+ tvjc = 0 tvje = 0 tvjs = 0
+ tis1 = 0 tise1 = 0 tisc1 = 0
+ tnf1 = -6e-3 tnr1 = 0 tne1 = 0 tnc1 = 0
+ tbf1 = 0 tbr1 = 0 tiss1 = 0 tvaf1 = 0
+ tvar1 = 0 tikf1 = 0 tikr1 = 0 tns1 = 0
+ trb1 = 0 trc1 = 0 tre1 = -0.005 tirb1 = 0
+ tsky130_fd_pr__res_generic_m1 = 0 tmjc1 = 0 tmje1 = 0 tmjs1 = 0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 0
+ tise2 = 0 tisc2 = 0 tnf2 = 0 tnr2 = 0
+ tne2 = 0 tnc2 = 0 tbf2 = 0 tbr2 = 0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 0
+ tikr2 = 0 tns2 = 0 trb2 = 0 trc2 = 0
+ tre2 = 0 tirb2 = 0 tsky130_fd_pr__res_generic_m2 = 0 tmjc2 = 0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0 titf2 = 0
+ ttr2 = 0
**************************************************************
*               QUASI
**************************************************************

.ends sky130_fd_pr__npn_11v0_W1p00L1p00
******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/02/23  UZMN (Usman Suriono)
*      Why     : New infrastructure of an npn model
*      What    : Converted from nsky130_fd_pr__pnp_05v5_W0p68L0p68ar1x2 model
*                Replaced all junction capacitance variation by correlated diodes.


.subckt  sky130_fd_pr__npn_05v5_W1p00L2p00 c b e s mult=1

+
+ 
.param  dkisnpn1x2 = 9.0950e-01
+ dkbfnpn1x2 = 9.6759e-01
+ var_is = {1/sw_func_rdn**2*(1+1.2*sw_mm_npn_is*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}
+ var_bf = {(sw_func_pw_rs*sw_pw_rs_mc)**2.2*(1+0.93*sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))}


Qsky130_fd_pr__npn_05v5_W1p00L2p00 c b e s nsky130_fd_pr__pnp_05v5_W0p68L0p68ar1x2_model 



.model nsky130_fd_pr__pnp_05v5_W0p68L0p68ar1x2_model npn level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ dcap = 2
+ cjc = '1.60339e-014*sw_func_pw_dnw_cj'
+ cje = '10.30981e-015*sw_func_nsd_pw_cj'
+ cjs = '3.05951e-014*sw_func_dnw_sub_cj'
+ fc = 0.5 mjc = 0.33982 mje = 0.44
+ mjs = 0.49 vjc = 0.58758 vje = 0.729 vjs = 0.5348
+ xcjc = 1 itf = '2.6e-03+7e-3' ptf = 20
+ tf = '6.34041e-011+4.5e-11'
+ tr = 0 vtf = '0.5+0.0' xtf = '2.0+0.9'
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.595 kf = 3.5568689e-11
**************************************************************
*               DC PARAMETERS
**************************************************************
+ is = '7.98e-018*dkisnpn1x2*var_is'
+ bf = '37.54*dkbfnpn1x2*var_bf'
+ vaf = '100 / var_bf'
+ ise = '5.77e-016*(1-sw_mm_npn_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult))'
+ nf = 1.0405 ikf = 0.0011462
+ subs = 1 rb = 885.61
+ re = 15.0 irb = 4.424e-005 rc = 61.677 rbm = 256.08
+ ne = 1.7924 ns = 1.0 br = 1
+ ibc = 0 iss = 0 nr = 0.96012
+ var = 0 ikr = 4.032e-008 nkf = 0.5 isc = 0
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xtb = 0 xti = 1.0713 eg = 1.188 gap1 = 0
+ gap2 = 0 ctc = 0
+ cte = 0 cts = 0 tlev = 0 tlevc = 0
+ tvjc = 0 tvje = 0 tvjs = 0
+ tis1 = 0 tise1 = 0 tisc1 = 0
+ tnf1 = 4.208e-005 tnr1 = -0.000522 tne1 = 0 tnc1 = 0
+ tbf1 = 0.00776 tbr1 = 0 tiss1 = 0 tvaf1 = 0
+ tvar1 = 0 tikf1 = -0.0074 tikr1 = 0 tns1 = 0
+ trb1 = 0 trc1 = 0 tre1 = 0 tirb1 = 0
+ tsky130_fd_pr__res_generic_m1 = 0 tmjc1 = 0 tmje1 = 0 tmjs1 = 0
+ ttf1 = 0 titf1 = 0 ttr1 = 0 tis2 = 4e-012
+ tise2 = 0 tisc2 = 0 tnf2 = -3.372e-007 tnr2 = 1.8e-006
+ tne2 = 0 tnc2 = 0 tbf2 = 6.48e-006 tbr2 = 0
+ tiss2 = 0 tvaf2 = 0 tvar2 = 0 tikf2 = 4e-005
+ tikr2 = 0 tns2 = 0 trb2 = 0 trc2 = 0
+ tre2 = 0 tirb2 = 0 tsky130_fd_pr__res_generic_m2 = 0 tmjc2 = 0
+ tmje2 = 0 tmjs2 = 0 ttf2 = 0 titf2 = 0
**************************************************************
*               QUASI
**************************************************************

.ends sky130_fd_pr__npn_05v5_W1p00L2p00
******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/02/19  UZMN (Usman Suriono)
*      Why     : New infrastructure of the sky130_fd_pr__pnp_05v5_W0p68L0p68 model
*      What    : Converted from sky130_fd_pr__pnp_05v5_W0p68L0p68par model
*                Changed the B-C capacitance variation from Pwell-Deep Nwell to
*                Nwell-Pwell (Nwell-Substrate cap is dominated by Nwell).
* Modified 03/08/2024  Tim Edwards  Removed substrate pin for backwards compatibility

.subckt  sky130_fd_pr__pnp_05v5_W3p40L3p40 c b e mult=1

+
+ 
.param  dkispp5x = 1.0046e+00
+ dkbfpp5x = 1.1288e+00
+ dknfpp5x = 1.0009e+00
+ dkisepp5x = 0.745
+ mm_bf = {0.45*sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult)}
+ mm_is = {0.13*sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_is*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult)}


Qsky130_fd_pr__pnp_05v5_W3p40L3p40 c b e c sky130_fd_pr__pnp_05v5_W0p68L0p68par5x_model 



.model sky130_fd_pr__pnp_05v5_W0p68L0p68par5x_model pnp level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30 subs = 1
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ cjc = '(9.155e-17*5.17*5.17+5.822e-16*4*5.17)*sw_func_nw_pw_cj'
+ cje = '(7.4079e-16*3.4*3.4+9.88e-17*4*3.4)*sw_func_psd_nw_cj'
+ cjs = 0
+ fc = 0.5 mjc = 0.24 mje = 0.3 mjs = 0.24
+ vjc = 0.54 vje = 0.74 vjs = 0.54 xcjc = 1
+ ptf = 0 tf = 6.15385e-010 tr = 5e-008 vtf = 1e-012
+ xtf = 0
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.30180 kf = 4.9435066e-011
**************************************************************
*               DC PARAMETERS
**************************************************************
+ bf = '16.603*dkbfpp5x*sw_nw_rs_mult**0.95*(1+mm_bf)'
+ ise = '1.0310e-015*dkisepp5x*(1-mm_bf)'
+ is = '7.1190e-018*dkispp5x / sw_func_rdp*(1+mm_is)'
+ vaf = '111.6 / sw_nw_rs_mult*(1-mm_bf)'
+ nf = '1.000*dknfpp5x'
+ rb = 73.32
+ re = 5.3848 irb = 0.0002
+ rc = 100.0 rbm = 25.19
+ ikf = 0.00038589 ne = 1.64
+ ns = 1 br = 0.2675 iss = 0 nr = 1
+ var = 4.3 ikr = 0.0043 nkf = 0.426 isc = 1.9855e-015
+ nc = 1.000
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xti = '5.0*( 1+mm_is)'
+ xtb = 1.692
+ eg = 1.125 tnf1 = 5.972e-006
+ tikf1 = -0.002456 tnf2 = -3.0e-008
**************************************************************
*               QUASI
**************************************************************

.ends sky130_fd_pr__pnp_05v5_W3p40L3p40
******************************************************************
******************************************************************
* *************************** Isolated Pwell Resistors ************************
* 2021/02/19  UZMN (Usman Suriono)
*      Why     : New infrastructure of the sky130_fd_pr__pnp_05v5_W0p68L0p68 model
*      What    : Converted from sky130_fd_pr__pnp_05v5_W0p68L0p68par model
* Modified 03/08/2024  Tim Edwards  Removed substrate pin for backwards compatibility

.subckt  sky130_fd_pr__pnp_05v5_W0p68L0p68 c b e mult=1

+
+ 
.param  dkbfpp = 9.5154e-01
+ dkispp = 9.2840e-01
+ mm_bf = {sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_bf*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult)}
+ mm_is = {sw_mm_sky130_fd_pr__pnp_05v5_W0p68L0p68_is*mismatch_factor*MC_MM_SWITCH*AGAUSS(0,1.0,1)/sqrt(mult)}

Qsky130_fd_pr__pnp_05v5_W0p68L0p68 c b e c sky130_fd_pr__pnp_05v5_W0p68L0p68_model 


**

.model sky130_fd_pr__pnp_05v5_W0p68L0p68_model pnp level = 1
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+ tref = 30
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+ cjc = 6.255e-015 cje = 6.113e-016 cjs = 0
+ fc = 0.5 mjc = 0.24 mje = 0.3 mjs = 0.24
+ vjc = 0.54 vje = 0.74 vjs = 0.54 xcjc = 1
+ ptf = 0 tf = 6.15385e-010 tr = 5e-008 vtf = 1e-12
+ xtf = 0
**************************************************************
*               Noise PARAMETERS
**************************************************************
+ af = 1.60722 kf = 4.9435066E-11
**************************************************************
*               DC PARAMETERS
**************************************************************
*+bf      = '19.35  * dkbfpp * (1 + 0.7*(sw_nw_rs_mult-1))   * (1 + mm_bf)'
+ bf = '19.35*dkbfpp*sw_nw_rs_mult**0.75*(1+mm_bf)'
+ ise = '9.4936e-017*(1-mm_bf)'
+ is = '1.5075e-018*dkispp / sw_func_rdp*(1+mm_is)'
+ vaf = '152.06 / sw_nw_rs_mult*(1-mm_bf)'
+ ikf = 3.3057e-005
+ rb = 316.21 re = 219 irb = 0.027411
+ rc = 531 rbm = 243.58
+ nf = '1.028'
+ ne = 1.6444
+ ns = 1 br = 0.2675 iss = 0 nr = 1
+ var = 4.3 ikr = 0.00043 nkf = 0.5 isc = 1.2e-015
+ nc = 1.003
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+ xti = {1.1*(1+mm_is)}
+ xtb = 2.2132 eg = 1.2 tikf1 = -0.0037823
+ tnf1 = 1.972e-006 tnf2 = -8.8e-007
**************************************************************
*               QUASI
**************************************************************

.ends sky130_fd_pr__pnp_05v5_W0p68L0p68

