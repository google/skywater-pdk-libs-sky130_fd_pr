* Copyright 2022 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SKY130 Spice File.
* Critical Model Parameters:
.param cnwvc = 0.0 + MC_PR_SWITCH*AGAUSS(0,1.0,1)

.param special_nfet_pass_lvt = 0.0 + MC_PR_SWITCH*AGAUSS(0,1.0,1)
* statistics {
*  process {
*     vary cnwvc dist=gauss std=1.0
*     vary special_nfet_pass_lvt dist=gauss std=1.0
*   }
*   mismatch {
*   }
* }
