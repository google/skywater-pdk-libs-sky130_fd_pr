# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__dfl1sd__example_168835116
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__dfl1sd__example_168835116 ;
  ORIGIN  0.180000  0.180000 ;
  SIZE  0.625000 BY  5.360000 ;
  OBS
    LAYER li1 ;
      RECT 0.055000 -0.020000 0.225000 4.730000 ;
  END
END sky130_fd_pr__dfl1sd__example_168835116
END LIBRARY
