# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__rf_sh_auvia__example_182061100
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__rf_sh_auvia__example_182061100 ;
  ORIGIN  4.710000  2.310000 ;
  SIZE  9.420000 BY  4.620000 ;
  OBS
    LAYER met4 ;
      RECT -4.710000 -2.310000 4.710000 2.310000 ;
    LAYER met5 ;
      RECT -4.710000 -2.310000 4.710000 2.310000 ;
    LAYER via4 ;
      RECT -4.590000 -2.190000 4.590000 2.190000 ;
  END
END sky130_fd_pr__rf_sh_auvia__example_182061100
END LIBRARY
