* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_nfet_01v8__toxe_slope=3.443e-03
.param sky130_fd_pr__special_nfet_01v8__lint_slope=0.0
.param sky130_fd_pr__special_nfet_01v8__nfactor_slope=0.0
.param sky130_fd_pr__special_nfet_01v8__voff_slope=0.007
.param sky130_fd_pr__special_nfet_01v8__vth0_slope=3.356e-03
.param sky130_fd_pr__special_nfet_01v8__vth0_slope1=7.356e-03
.param sky130_fd_pr__special_nfet_01v8__wint_slope=0
